VERSION	5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    CAPACITANCE PICOFARADS 10 ;
    CURRENT MILLIAMPS 10000 ;
    VOLTAGE VOLTS 1000 ;
    DATABASE MICRONS 2000 ;
END UNITS
MANUFACTURINGGRID 0.005 ;
LAYER PO
    TYPE MASTERSLICE ;
END PO
LAYER CO
    TYPE CUT ;
END CO
LAYER M1
    TYPE ROUTING ;
    DIRECTION	HORIZONTAL ;
    PITCH	0.140 ;
    OFFSET	0.000 ;
    HEIGHT	0.53500 ;
    THICKNESS	0.12500 ;
    WIDTH	0.070 ;
    SPACING 0.070 ;
    AREA	0.0215 ;
 
	
    RESISTANCE RPERSQ 0.3080000000 ;
    CAPACITANCE CPERSQDIST 0.0002317460 ;
    EDGECAPACITANCE	0.0000808000 ;
END M1
LAYER VIA1
    TYPE CUT ;
    SPACING	0.095 ;
END VIA1
LAYER M2
    TYPE ROUTING ;
    DIRECTION	VERTICAL ;
    PITCH	0.140 ;
    OFFSET	0.070 ;
    HEIGHT	0.78000 ;
    THICKNESS	0.14000 ;
    WIDTH	0.070 ;
    SPACING 0.070 ;
    AREA	0.027 ;
 
  
    RESISTANCE RPERSQ 0.2780000000 ;
    CAPACITANCE CPERSQDIST 0.0003444444 ;
    EDGECAPACITANCE	0.0000730000 ;
END M2
LAYER VIA2
    TYPE CUT ;
    SPACING	0.095 ;
END VIA2
LAYER M3
    TYPE ROUTING ;
    DIRECTION	HORIZONTAL ;
    PITCH	0.140 ;
    OFFSET	0.000 ;
    HEIGHT	1.04000 ;
    THICKNESS	0.14000 ;
    WIDTH	0.070 ;
    SPACING 0.070 ;
    AREA	0.027 ;
 
  
    RESISTANCE RPERSQ 0.2780000000 ;
    CAPACITANCE CPERSQDIST 0.0003444444 ;
    EDGECAPACITANCE	0.0000730000 ;
END M3
LAYER VIA3
    TYPE CUT ;
    SPACING	0.095 ;
END VIA3
LAYER M4
    TYPE ROUTING ;
    DIRECTION	VERTICAL ;
    PITCH	0.140 ;
    OFFSET	0.070 ;
    HEIGHT	1.30000 ;
    THICKNESS	0.14000 ;
    WIDTH	0.070 ;
    SPACING 0.070 ;
    AREA	0.027 ;
 
  
  
    RESISTANCE RPERSQ 0.2780000000 ;
    CAPACITANCE CPERSQDIST 0.0003444444 ;
    EDGECAPACITANCE	0.0000730000 ;
END M4
LAYER VIA4
    TYPE CUT ;
    SPACING	0.095 ;
END VIA4
LAYER M5
    TYPE ROUTING ;
    DIRECTION	HORIZONTAL ;
    PITCH	0.140 ;
    OFFSET	0.000 ;
    HEIGHT	1.56000 ;
    THICKNESS	0.14000 ;
    WIDTH	0.070 ;
    SPACING 0.070 ;
    AREA	0.027 ;
 
  
  
    RESISTANCE RPERSQ 0.2780000000 ;
    CAPACITANCE CPERSQDIST 0.0003444444 ;
    EDGECAPACITANCE	0.0000730000 ;
END M5
LAYER VIA5
    TYPE CUT ;
    SPACING	0.095 ;
END VIA5
LAYER M6
    TYPE ROUTING ;
    DIRECTION	VERTICAL ;
    PITCH	0.140 ;
    OFFSET	0.070 ;
    HEIGHT	1.82000 ;
    THICKNESS	0.14000 ;
    WIDTH	0.070 ;
    SPACING 0.070 ;
    AREA	0.027 ;
 
  
  
    RESISTANCE RPERSQ 0.2780000000 ;
    CAPACITANCE CPERSQDIST 0.0003444444 ;
    EDGECAPACITANCE	0.0000730000 ;
END M6
LAYER VIA6
    TYPE CUT ;
    SPACING	0.340 ;
END VIA6
LAYER M7
    TYPE ROUTING ;
    DIRECTION	HORIZONTAL ;
    PITCH	0.800 ;
    OFFSET	0.000 ;
    HEIGHT	2.55500 ;
    THICKNESS	0.85000 ;
    WIDTH	0.400 ;
    SPACING 0.400 ;
    AREA	0.565 ;
  
    RESISTANCE RPERSQ 0.0220000000 ;
    CAPACITANCE CPERSQDIST 0.0000613889 ;
    EDGECAPACITANCE	0.0000912000 ;
END M7
LAYER VIA7
    TYPE CUT ;
    SPACING	0.340 ;
END VIA7
LAYER M8
    TYPE ROUTING ;
    DIRECTION	VERTICAL ;
    PITCH	0.800 ;
    OFFSET	0.070 ;
    HEIGHT	4.00000 ;
    THICKNESS	0.85000 ;
    WIDTH	0.400 ;
    SPACING 0.400 ;
    AREA	0.565 ;
  
    RESISTANCE RPERSQ 0.0220000000 ;
    CAPACITANCE CPERSQDIST 0.0000613889 ;
    EDGECAPACITANCE	0.0000935000 ;
END M8
LAYER OVERLAP
    TYPE OVERLAP ;
END OVERLAP
VIA VIA12_1cut DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M1 ;
        RECT -0.065 -0.035  0.065  0.035 ;
    LAYER VIA1 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M2 ;
        RECT -0.035 -0.065  0.035  0.065 ;
END VIA12_1cut
VIA VIA12_1cut_H DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M1 ;
        RECT -0.065 -0.035  0.065  0.035 ;
    LAYER VIA1 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M2 ;
        RECT -0.065 -0.035  0.065  0.035 ;
END VIA12_1cut_H
                 
VIA VIA12_1cut_V DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M1 ;
        RECT -0.035 -0.065  0.035  0.065 ;
    LAYER VIA1 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M2 ;
        RECT -0.035 -0.065  0.035  0.065 ;
END VIA12_1cut_V
VIA VIA12_1cut_FAT_C DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M1 ;
        RECT -0.085 -0.035  0.085  0.035 ;
    LAYER VIA1 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M2 ;
        RECT -0.035 -0.085  0.035  0.085 ;
END VIA12_1cut_FAT_C
             
VIA VIA12_1cut_FAT_H DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M1 ;
        RECT -0.085 -0.035  0.085  0.035 ;
    LAYER VIA1 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M2 ;
        RECT -0.085 -0.035  0.085  0.035 ;
END VIA12_1cut_FAT_H
VIA VIA12_1cut_FAT_V DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M1 ;
        RECT -0.035 -0.085  0.035  0.085 ;
    LAYER VIA1 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M2 ;
        RECT -0.035 -0.085  0.035  0.085 ;
END VIA12_1cut_FAT_V
VIA VIA12_1cut_FAT DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M1 ;
        RECT -0.065 -0.065  0.065  0.065 ;
    LAYER VIA1 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M2 ;
        RECT -0.065 -0.065  0.065  0.065 ;
END VIA12_1cut_FAT
                 
VIA VIA12_1cut_R90 DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M1 ;
        RECT -0.035 -0.065  0.035  0.065 ;
    LAYER VIA1 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M2 ;
        RECT -0.065 -0.035  0.065  0.035 ;
END VIA12_1cut_R90
VIA VIA12_2cut_E DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M1 ;
        RECT -0.065 -0.035  0.205  0.035 ;
    LAYER VIA1 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT 0.105 -0.035  0.175  0.035 ;
    LAYER M2 ;
        RECT -0.035 -0.065  0.175  0.065 ;
END VIA12_2cut_E
VIA VIA12_2cut_E_FB DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M1 ;
       RECT -0.065 -0.065 0.205 0.065 ;
    LAYER VIA1 ;
        RECT -0.035 -0.035 0.035 0.035 ;
        RECT 0.105 -0.035 0.175 0.035 ;
    LAYER M2 ;
       RECT -0.065 -0.065 0.205 0.065 ;
END VIA12_2cut_E_FB
VIA VIA12_2cut_W DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M1 ;
        RECT -0.205 -0.035  0.065  0.035 ;
    LAYER VIA1 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT -0.175 -0.035  -0.105  0.035 ;
    LAYER M2 ;
        RECT -0.175 -0.065  0.035  0.065 ;
END VIA12_2cut_W
VIA VIA12_2cut_W_FB DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M1 ;
       RECT -0.205 -0.065 0.065 0.065 ;
    LAYER VIA1 ;
        RECT -0.035 -0.035 0.035 0.035 ;
        RECT -0.175 -0.035 -0.105 0.035 ;
    LAYER M2 ;
       RECT -0.205 -0.065 0.065 0.065 ;
END VIA12_2cut_W_FB
VIA VIA12_2cut_N DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M1 ;
        RECT -0.065 -0.035  0.065  0.175 ;
    LAYER VIA1 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT -0.035 0.105  0.035  0.175 ;
    LAYER M2 ;
        RECT -0.035 -0.065  0.035  0.205 ;
END VIA12_2cut_N
VIA VIA12_2cut_N_FB DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M1 ;
       RECT -0.065 -0.065 0.065 0.205 ;
    LAYER VIA1 ;
        RECT -0.035 -0.035 0.035 0.035 ;
        RECT -0.035 0.105 0.035 0.175 ;
    LAYER M2 ;
       RECT -0.065 -0.065 0.065 0.205 ;
END VIA12_2cut_N_FB
VIA VIA12_2cut_S DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M1 ;
        RECT -0.065 -0.175  0.065  0.035 ;
    LAYER VIA1 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT -0.035 -0.175  0.035  -0.105 ;
    LAYER M2 ;
        RECT -0.035 -0.205  0.035  0.065 ;
END VIA12_2cut_S
VIA VIA12_2cut_S_FB DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M1 ;
       RECT -0.065 -0.205 0.065 0.065 ;
    LAYER VIA1 ;
        RECT -0.035 -0.035 0.035 0.035 ;
        RECT -0.035 -0.175 0.035 -0.105 ;
    LAYER M2 ;
       RECT -0.065 -0.205 0.065 0.065 ;
END VIA12_2cut_S_FB
VIA VIA12_2cut_HN DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M1 ;
        RECT -0.035 -0.065  0.035  0.235 ;
    LAYER VIA1 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT -0.035 0.135  0.035  0.205 ;
    LAYER M2 ;
        RECT -0.035 -0.065  0.035  0.235 ;
END VIA12_2cut_HN
 
VIA VIA12_2cut_HS DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M1 ;
        RECT -0.035 -0.235  0.035  0.065 ;
    LAYER VIA1 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT -0.035 -0.205  0.035  -0.135 ;
    LAYER M2 ;
        RECT -0.035 -0.235  0.035  0.065 ;
END VIA12_2cut_HS
VIA VIA12_4cut DEFAULT
    RESISTANCE 1.6750000000 ;
    LAYER M1 ;
        RECT -0.135 -0.105  0.135  0.105 ;
    LAYER VIA1 ;
        RECT -0.105 -0.105  -0.035  -0.035 ;
        RECT -0.105 0.035  -0.035  0.105 ;
        RECT 0.035 0.035  0.105  0.105 ;
        RECT 0.035 -0.105  0.105  -0.035 ;
    LAYER M2 ;
        RECT -0.105 -0.135  0.105  0.135 ;
END VIA12_4cut
VIA VIA23_1cut DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M2 ;
        RECT -0.035 -0.065  0.035  0.065 ;
    LAYER VIA2 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M3 ;
        RECT -0.065 -0.035  0.065  0.035 ;
END VIA23_1cut
VIA VIA23_1cut_V DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M2 ;
        RECT -0.035 -0.065  0.035  0.065 ;
    LAYER VIA2 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M3 ;
        RECT -0.035 -0.065  0.035  0.065 ;
END VIA23_1cut_V
VIA VIA23_1cut_H DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M2 ;
        RECT -0.065 -0.035  0.065  0.035 ;
    LAYER VIA2 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M3 ;
        RECT -0.065 -0.035  0.065  0.035 ;
END VIA23_1cut_H
VIA VIA23_1cut_FAT_C DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M2 ;
        RECT -0.035 -0.085  0.035  0.085 ;
    LAYER VIA2 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M3 ;
        RECT -0.085 -0.035  0.085  0.035 ;
END VIA23_1cut_FAT_C
             
VIA VIA23_1cut_FAT_V DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M2 ;
        RECT -0.035 -0.085  0.035  0.085 ;
    LAYER VIA2 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M3 ;
        RECT -0.035 -0.085  0.035  0.085 ;
END VIA23_1cut_FAT_V
VIA VIA23_1cut_FAT_H DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M2 ;
        RECT -0.085 -0.035  0.085  0.035 ;
    LAYER VIA2 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M3 ;
        RECT -0.085 -0.035  0.085  0.035 ;
END VIA23_1cut_FAT_H
VIA VIA23_1cut_FAT DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M2 ;
        RECT -0.065 -0.065  0.065  0.065 ;
    LAYER VIA2 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M3 ;
        RECT -0.065 -0.065  0.065  0.065 ;
END VIA23_1cut_FAT
                 
VIA VIA23_1stack_N DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M2 ;
        RECT -0.035 -0.065  0.035  0.325 ;
    LAYER VIA2 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M3 ;
        RECT -0.065 -0.035  0.065  0.035 ;
END VIA23_1stack_N
VIA VIA23_1stack_S DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M2 ;
        RECT -0.035 -0.325  0.035  0.065 ;
    LAYER VIA2 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M3 ;
        RECT -0.065 -0.035  0.065  0.035 ;
END VIA23_1stack_S
VIA VIA23_2cut_E DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M2 ;
        RECT -0.035 -0.065  0.175  0.065 ;
    LAYER VIA2 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT 0.105 -0.035  0.175  0.035 ;
    LAYER M3 ;
        RECT -0.065 -0.035  0.205  0.035 ;
END VIA23_2cut_E
VIA VIA23_2cut_E_FB DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M2 ;
       RECT -0.065 -0.065 0.205 0.065 ;
    LAYER VIA2 ;
        RECT -0.035 -0.035 0.035 0.035 ;
        RECT 0.105 -0.035 0.175 0.035 ;
    LAYER M3 ;
       RECT -0.065 -0.065 0.205 0.065 ;
END VIA23_2cut_E_FB
 
VIA VIA23_2cut_W DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M2 ;
        RECT -0.175 -0.065  0.035  0.065 ;
    LAYER VIA2 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT -0.175 -0.035  -0.105  0.035 ;
    LAYER M3 ;
        RECT -0.205 -0.035  0.065  0.035 ;
END VIA23_2cut_W
VIA VIA23_2cut_W_FB DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M2 ;
       RECT -0.205 -0.065 0.065 0.065 ;
    LAYER VIA2 ;
        RECT -0.035 -0.035 0.035 0.035 ;
        RECT -0.175 -0.035 -0.105 0.035 ;
    LAYER M3 ;
       RECT -0.205 -0.065 0.065 0.065 ;
END VIA23_2cut_W_FB
 
VIA VIA23_2cut_N DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M2 ;
        RECT -0.035 -0.065  0.035  0.205 ;
    LAYER VIA2 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT -0.035 0.105  0.035  0.175 ;
    LAYER M3 ;
        RECT -0.065 -0.035  0.065  0.175 ;
END VIA23_2cut_N
VIA VIA23_2cut_N_FB DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M2 ;
       RECT -0.065 -0.065 0.065 0.205 ;
    LAYER VIA2 ;
        RECT -0.035 -0.035 0.035 0.035 ;
        RECT -0.035 0.105 0.035 0.175 ;
    LAYER M3 ;
       RECT -0.065 -0.065 0.065 0.205 ;
END VIA23_2cut_N_FB
 
VIA VIA23_2cut_S DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M2 ;
        RECT -0.035 -0.205  0.035  0.065 ;
    LAYER VIA2 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT -0.035 -0.175  0.035  -0.105 ;
    LAYER M3 ;
        RECT -0.065 -0.175  0.065  0.035 ;
END VIA23_2cut_S
VIA VIA23_2cut_S_FB DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M2 ;
       RECT -0.065 -0.205 0.065 0.065 ;
    LAYER VIA2 ;
        RECT -0.035 -0.035 0.035 0.035 ;
        RECT -0.035 -0.175 0.035 -0.105 ;
    LAYER M3 ;
       RECT -0.065 -0.205 0.065 0.065 ;
END VIA23_2cut_S_FB
VIA VIA23_4cut DEFAULT
    RESISTANCE 1.6750000000 ;
    LAYER M2 ;
        RECT -0.105 -0.135  0.105  0.135 ;
    LAYER VIA2 ;
        RECT -0.105 -0.105  -0.035  -0.035 ;
        RECT -0.105 0.035  -0.035  0.105 ;
        RECT 0.035 0.035  0.105  0.105 ;
        RECT 0.035 -0.105  0.105  -0.035 ;
    LAYER M3 ;
        RECT -0.135 -0.105  0.135  0.105 ;
END VIA23_4cut
VIA VIA34_1cut DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M3 ;
        RECT -0.065 -0.035  0.065  0.035 ;
    LAYER VIA3 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M4 ;
        RECT -0.035 -0.065  0.035  0.065 ;
END VIA34_1cut
VIA VIA34_1cut_H DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M3 ;
        RECT -0.065 -0.035  0.065  0.035 ;
    LAYER VIA3 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M4 ;
        RECT -0.065 -0.035  0.065  0.035 ;
END VIA34_1cut_H
                 
VIA VIA34_1cut_V DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M3 ;
        RECT -0.035 -0.065  0.035  0.065 ;
    LAYER VIA3 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M4 ;
        RECT -0.035 -0.065  0.035  0.065 ;
END VIA34_1cut_V
VIA VIA34_1cut_FAT_C DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M3 ;
        RECT -0.085 -0.035  0.085  0.035 ;
    LAYER VIA3 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M4 ;
        RECT -0.035 -0.085  0.035  0.085 ;
END VIA34_1cut_FAT_C
             
VIA VIA34_1cut_FAT_H DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M3 ;
        RECT -0.085 -0.035  0.085  0.035 ;
    LAYER VIA3 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M4 ;
        RECT -0.085 -0.035  0.085  0.035 ;
END VIA34_1cut_FAT_H
VIA VIA34_1cut_FAT_V DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M3 ;
        RECT -0.035 -0.085  0.035  0.085 ;
    LAYER VIA3 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M4 ;
        RECT -0.035 -0.085  0.035  0.085 ;
END VIA34_1cut_FAT_V
VIA VIA34_1cut_FAT DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M3 ;
        RECT -0.065 -0.065  0.065  0.065 ;
    LAYER VIA3 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M4 ;
        RECT -0.065 -0.065  0.065  0.065 ;
END VIA34_1cut_FAT
                 
VIA VIA34_1stack_E DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M3 ;
        RECT -0.065 -0.035  0.325  0.035 ;
    LAYER VIA3 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M4 ;
        RECT -0.035 -0.065  0.035  0.065 ;
END VIA34_1stack_E
VIA VIA34_1stack_W DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M3 ;
        RECT -0.325 -0.035  0.065  0.035 ;
    LAYER VIA3 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M4 ;
        RECT -0.035 -0.065  0.035  0.065 ;
END VIA34_1stack_W
VIA VIA34_2cut_E DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M3 ;
        RECT -0.065 -0.035  0.205  0.035 ;
    LAYER VIA3 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT 0.105 -0.035  0.175  0.035 ;
    LAYER M4 ;
        RECT -0.035 -0.065  0.175  0.065 ;
END VIA34_2cut_E
VIA VIA34_2cut_E_FB DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M3 ;
       RECT -0.065 -0.065 0.205 0.065 ;
    LAYER VIA3 ;
        RECT -0.035 -0.035 0.035 0.035 ;
        RECT 0.105 -0.035 0.175 0.035 ;
    LAYER M4 ;
       RECT -0.065 -0.065 0.205 0.065 ;
END VIA34_2cut_E_FB
 
VIA VIA34_2cut_W DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M3 ;
        RECT -0.205 -0.035  0.065  0.035 ;
    LAYER VIA3 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT -0.175 -0.035  -0.105  0.035 ;
    LAYER M4 ;
        RECT -0.175 -0.065  0.035  0.065 ;
END VIA34_2cut_W
VIA VIA34_2cut_W_FB DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M3 ;
       RECT -0.205 -0.065 0.065 0.065 ;
    LAYER VIA3 ;
        RECT -0.035 -0.035 0.035 0.035 ;
        RECT -0.175 -0.035 -0.105 0.035 ;
    LAYER M4 ;
       RECT -0.205 -0.065 0.065 0.065 ;
END VIA34_2cut_W_FB
 
VIA VIA34_2cut_N DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M3 ;
        RECT -0.065 -0.035  0.065  0.175 ;
    LAYER VIA3 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT -0.035 0.105  0.035  0.175 ;
    LAYER M4 ;
        RECT -0.035 -0.065  0.035  0.205 ;
END VIA34_2cut_N
VIA VIA34_2cut_N_FB DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M3 ;
       RECT -0.065 -0.065 0.065 0.205 ;
    LAYER VIA3 ;
        RECT -0.035 -0.035 0.035 0.035 ;
        RECT -0.035 0.105 0.035 0.175 ;
    LAYER M4 ;
       RECT -0.065 -0.065 0.065 0.205 ;
END VIA34_2cut_N_FB
 
VIA VIA34_2cut_S DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M3 ;
        RECT -0.065 -0.175  0.065  0.035 ;
    LAYER VIA3 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT -0.035 -0.175  0.035  -0.105 ;
    LAYER M4 ;
        RECT -0.035 -0.205  0.035  0.065 ;
END VIA34_2cut_S
VIA VIA34_2cut_S_FB DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M3 ;
       RECT -0.065 -0.205 0.065 0.065 ;
    LAYER VIA3 ;
        RECT -0.035 -0.035 0.035 0.035 ;
        RECT -0.035 -0.175 0.035 -0.105 ;
    LAYER M4 ;
       RECT -0.065 -0.205 0.065 0.065 ;
END VIA34_2cut_S_FB
VIA VIA34_4cut DEFAULT
    RESISTANCE 1.6750000000 ;
    LAYER M3 ;
        RECT -0.135 -0.105  0.135  0.105 ;
    LAYER VIA3 ;
        RECT -0.105 -0.105  -0.035  -0.035 ;
        RECT -0.105 0.035  -0.035  0.105 ;
        RECT 0.035 0.035  0.105  0.105 ;
        RECT 0.035 -0.105  0.105  -0.035 ;
    LAYER M4 ;
        RECT -0.105 -0.135  0.105  0.135 ;
END VIA34_4cut
VIA VIA45_1cut DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M4 ;
        RECT -0.035 -0.065  0.035  0.065 ;
    LAYER VIA4 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M5 ;
        RECT -0.065 -0.035  0.065  0.035 ;
END VIA45_1cut
VIA VIA45_1cut_V DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M4 ;
        RECT -0.035 -0.065  0.035  0.065 ;
    LAYER VIA4 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M5 ;
        RECT -0.035 -0.065  0.035  0.065 ;
END VIA45_1cut_V
VIA VIA45_1cut_H DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M4 ;
        RECT -0.065 -0.035  0.065  0.035 ;
    LAYER VIA4 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M5 ;
        RECT -0.065 -0.035  0.065  0.035 ;
END VIA45_1cut_H
VIA VIA45_1cut_FAT_C DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M4 ;
        RECT -0.035 -0.085  0.035  0.085 ;
    LAYER VIA4 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M5 ;
        RECT -0.085 -0.035  0.085  0.035 ;
END VIA45_1cut_FAT_C
             
VIA VIA45_1cut_FAT_V DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M4 ;
        RECT -0.035 -0.085  0.035  0.085 ;
    LAYER VIA4 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M5 ;
        RECT -0.035 -0.085  0.035  0.085 ;
END VIA45_1cut_FAT_V
VIA VIA45_1cut_FAT_H DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M4 ;
        RECT -0.085 -0.035  0.085  0.035 ;
    LAYER VIA4 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M5 ;
        RECT -0.085 -0.035  0.085  0.035 ;
END VIA45_1cut_FAT_H
VIA VIA45_1cut_FAT DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M4 ;
        RECT -0.065 -0.065  0.065  0.065 ;
    LAYER VIA4 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M5 ;
        RECT -0.065 -0.065  0.065  0.065 ;
END VIA45_1cut_FAT
                 
VIA VIA45_1stack_N DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M4 ;
        RECT -0.035 -0.065  0.035  0.325 ;
    LAYER VIA4 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M5 ;
        RECT -0.065 -0.035  0.065  0.035 ;
END VIA45_1stack_N
VIA VIA45_1stack_S DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M4 ;
        RECT -0.035 -0.325  0.035  0.065 ;
    LAYER VIA4 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M5 ;
        RECT -0.065 -0.035  0.065  0.035 ;
END VIA45_1stack_S
VIA VIA45_2cut_E DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M4 ;
        RECT -0.035 -0.065  0.175  0.065 ;
    LAYER VIA4 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT 0.105 -0.035  0.175  0.035 ;
    LAYER M5 ;
        RECT -0.065 -0.035  0.205  0.035 ;
END VIA45_2cut_E
VIA VIA45_2cut_E_FB DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M4 ;
       RECT -0.065 -0.065 0.205 0.065 ;
    LAYER VIA4 ;
        RECT -0.035 -0.035 0.035 0.035 ;
        RECT 0.105 -0.035 0.175 0.035 ;
    LAYER M5 ;
       RECT -0.065 -0.065 0.205 0.065 ;
END VIA45_2cut_E_FB
 
VIA VIA45_2cut_W DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M4 ;
        RECT -0.175 -0.065  0.035  0.065 ;
    LAYER VIA4 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT -0.175 -0.035  -0.105  0.035 ;
    LAYER M5 ;
        RECT -0.205 -0.035  0.065  0.035 ;
END VIA45_2cut_W
VIA VIA45_2cut_W_FB DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M4 ;
       RECT -0.205 -0.065 0.065 0.065 ;
    LAYER VIA4 ;
        RECT -0.035 -0.035 0.035 0.035 ;
        RECT -0.175 -0.035 -0.105 0.035 ;
    LAYER M5 ;
       RECT -0.205 -0.065 0.065 0.065 ;
END VIA45_2cut_W_FB
 
VIA VIA45_2cut_N DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M4 ;
        RECT -0.035 -0.065  0.035  0.205 ;
    LAYER VIA4 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT -0.035 0.105  0.035  0.175 ;
    LAYER M5 ;
        RECT -0.065 -0.035  0.065  0.175 ;
END VIA45_2cut_N
VIA VIA45_2cut_N_FB DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M4 ;
       RECT -0.065 -0.065 0.065 0.205 ;
    LAYER VIA4 ;
        RECT -0.035 -0.035 0.035 0.035 ;
        RECT -0.035 0.105 0.035 0.175 ;
    LAYER M5 ;
       RECT -0.065 -0.065 0.065 0.205 ;
END VIA45_2cut_N_FB
 
VIA VIA45_2cut_S DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M4 ;
        RECT -0.035 -0.205  0.035  0.065 ;
    LAYER VIA4 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT -0.035 -0.175  0.035  -0.105 ;
    LAYER M5 ;
        RECT -0.065 -0.175  0.065  0.035 ;
END VIA45_2cut_S
VIA VIA45_2cut_S_FB DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M4 ;
       RECT -0.065 -0.205 0.065 0.065 ;
    LAYER VIA4 ;
        RECT -0.035 -0.035 0.035 0.035 ;
        RECT -0.035 -0.175 0.035 -0.105 ;
    LAYER M5 ;
       RECT -0.065 -0.205 0.065 0.065 ;
END VIA45_2cut_S_FB
VIA VIA45_4cut DEFAULT
    RESISTANCE 1.6750000000 ;
    LAYER M4 ;
        RECT -0.105 -0.135  0.105  0.135 ;
    LAYER VIA4 ;
        RECT -0.105 -0.105  -0.035  -0.035 ;
        RECT -0.105 0.035  -0.035  0.105 ;
        RECT 0.035 0.035  0.105  0.105 ;
        RECT 0.035 -0.105  0.105  -0.035 ;
    LAYER M5 ;
        RECT -0.135 -0.105  0.135  0.105 ;
END VIA45_4cut
VIA VIA56_1cut DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M5 ;
        RECT -0.065 -0.035  0.065  0.035 ;
    LAYER VIA5 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M6 ;
        RECT -0.035 -0.065  0.035  0.065 ;
END VIA56_1cut
VIA VIA56_1cut_H DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M5 ;
        RECT -0.065 -0.035  0.065  0.035 ;
    LAYER VIA5 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M6 ;
        RECT -0.065 -0.035  0.065  0.035 ;
END VIA56_1cut_H
                 
VIA VIA56_1cut_V DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M5 ;
        RECT -0.035 -0.065  0.035  0.065 ;
    LAYER VIA5 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M6 ;
        RECT -0.035 -0.065  0.035  0.065 ;
END VIA56_1cut_V
VIA VIA56_1cut_FAT_C DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M5 ;
        RECT -0.085 -0.035  0.085  0.035 ;
    LAYER VIA5 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M6 ;
        RECT -0.035 -0.085  0.035  0.085 ;
END VIA56_1cut_FAT_C
             
VIA VIA56_1cut_FAT_H DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M5 ;
        RECT -0.085 -0.035  0.085  0.035 ;
    LAYER VIA5 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M6 ;
        RECT -0.085 -0.035  0.085  0.035 ;
END VIA56_1cut_FAT_H
VIA VIA56_1cut_FAT_V DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M5 ;
        RECT -0.035 -0.085  0.035  0.085 ;
    LAYER VIA5 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M6 ;
        RECT -0.035 -0.085  0.035  0.085 ;
END VIA56_1cut_FAT_V
VIA VIA56_1cut_FAT DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M5 ;
        RECT -0.065 -0.065  0.065  0.065 ;
    LAYER VIA5 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M6 ;
        RECT -0.065 -0.065  0.065  0.065 ;
END VIA56_1cut_FAT
                 
VIA VIA56_1stack_E DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M5 ;
        RECT -0.065 -0.035  0.325  0.035 ;
    LAYER VIA5 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M6 ;
        RECT -0.035 -0.065  0.035  0.065 ;
END VIA56_1stack_E
VIA VIA56_1stack_W DEFAULT
    RESISTANCE 6.7000000000 ;
    LAYER M5 ;
        RECT -0.325 -0.035  0.065  0.035 ;
    LAYER VIA5 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M6 ;
        RECT -0.035 -0.065  0.035  0.065 ;
END VIA56_1stack_W
VIA VIA56_2cut_E DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M5 ;
        RECT -0.065 -0.035  0.205  0.035 ;
    LAYER VIA5 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT 0.105 -0.035  0.175  0.035 ;
    LAYER M6 ;
        RECT -0.035 -0.065  0.175  0.065 ;
END VIA56_2cut_E
VIA VIA56_2cut_E_FB DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M5 ;
       RECT -0.065 -0.065 0.205 0.065 ;
    LAYER VIA5 ;
        RECT -0.035 -0.035 0.035 0.035 ;
        RECT 0.105 -0.035 0.175 0.035 ;
    LAYER M6 ;
       RECT -0.065 -0.065 0.205 0.065 ;
END VIA56_2cut_E_FB
 
VIA VIA56_2cut_W DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M5 ;
        RECT -0.205 -0.035  0.065  0.035 ;
    LAYER VIA5 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT -0.175 -0.035  -0.105  0.035 ;
    LAYER M6 ;
        RECT -0.175 -0.065  0.035  0.065 ;
END VIA56_2cut_W
VIA VIA56_2cut_W_FB DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M5 ;
       RECT -0.205 -0.065 0.065 0.065 ;
    LAYER VIA5 ;
        RECT -0.035 -0.035 0.035 0.035 ;
        RECT -0.175 -0.035 -0.105 0.035 ;
    LAYER M6 ;
       RECT -0.205 -0.065 0.065 0.065 ;
END VIA56_2cut_W_FB
 
VIA VIA56_2cut_N DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M5 ;
        RECT -0.065 -0.035  0.065  0.175 ;
    LAYER VIA5 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT -0.035 0.105  0.035  0.175 ;
    LAYER M6 ;
        RECT -0.035 -0.065  0.035  0.205 ;
END VIA56_2cut_N
VIA VIA56_2cut_N_FB DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M5 ;
       RECT -0.065 -0.065 0.065 0.205 ;
    LAYER VIA5 ;
        RECT -0.035 -0.035 0.035 0.035 ;
        RECT -0.035 0.105 0.035 0.175 ;
    LAYER M6 ;
       RECT -0.065 -0.065 0.065 0.205 ;
END VIA56_2cut_N_FB
 
VIA VIA56_2cut_S DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M5 ;
        RECT -0.065 -0.175  0.065  0.035 ;
    LAYER VIA5 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT -0.035 -0.175  0.035  -0.105 ;
    LAYER M6 ;
        RECT -0.035 -0.205  0.035  0.065 ;
END VIA56_2cut_S
VIA VIA56_2cut_S_FB DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M5 ;
       RECT -0.065 -0.205 0.065 0.065 ;
    LAYER VIA5 ;
        RECT -0.035 -0.035 0.035 0.035 ;
        RECT -0.035 -0.175 0.035 -0.105 ;
    LAYER M6 ;
       RECT -0.065 -0.205 0.065 0.065 ;
END VIA56_2cut_S_FB
VIA VIA56_2stack_E DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M5 ;
        RECT -0.065 -0.035  0.325  0.035 ;
    LAYER VIA5 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT 0.105 -0.035  0.175  0.035 ;
    LAYER M6 ;
        RECT -0.035 -0.065  0.175  0.065 ;
END VIA56_2stack_E
 
VIA VIA56_2stack_W DEFAULT
    RESISTANCE 3.3500000000 ;
    LAYER M5 ;
        RECT -0.325 -0.035  0.065  0.035 ;
    LAYER VIA5 ;
        RECT -0.035 -0.035  0.035  0.035 ;
        RECT -0.175 -0.035  -0.105  0.035 ;
    LAYER M6 ;
        RECT -0.175 -0.065  0.035  0.065 ;
END VIA56_2stack_W
VIA VIA56_4cut DEFAULT
    RESISTANCE 1.6750000000 ;
    LAYER M5 ;
        RECT -0.135 -0.105  0.135  0.105 ;
    LAYER VIA5 ;
        RECT -0.105 -0.105  -0.035  -0.035 ;
        RECT -0.105 0.035  -0.035  0.105 ;
        RECT 0.035 0.035  0.105  0.105 ;
        RECT 0.035 -0.105  0.105  -0.035 ;
    LAYER M6 ;
        RECT -0.105 -0.135  0.105  0.135 ;
END VIA56_4cut
VIA VIA67_1cut DEFAULT
    RESISTANCE 0.2700000000 ;
    LAYER M6 ;
        RECT -0.200 -0.260  0.200  0.260 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.200 ;
END VIA67_1cut
VIA VIA67_1cut_H DEFAULT
    RESISTANCE 0.2700000000 ;
    LAYER M6 ;
        RECT -0.260 -0.200  0.260  0.200 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.200 ;
END VIA67_1cut_H
                 
VIA VIA67_1cut_V DEFAULT
    RESISTANCE 0.2700000000 ;
    LAYER M6 ;
        RECT -0.200 -0.260  0.200  0.260 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.200 -0.260  0.200  0.260 ;
END VIA67_1cut_V
VIA VIA67_1cut_FAT_C DEFAULT
    RESISTANCE 0.2700000000 ;
    LAYER M6 ;
        RECT -0.200 -0.260  0.200  0.260 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.200 ;
END VIA67_1cut_FAT_C
VIA VIA67_1cut_FAT_H DEFAULT
    RESISTANCE 0.2700000000 ;
    LAYER M6 ;
        RECT -0.260 -0.200  0.260  0.200 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.200 ;
END VIA67_1cut_FAT_H
VIA VIA67_1cut_FAT_V DEFAULT
    RESISTANCE 0.2700000000 ;
    LAYER M6 ;
        RECT -0.200 -0.260  0.200  0.260 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.200 -0.260  0.200  0.260 ;
END VIA67_1cut_FAT_V
VIA VIA67_1cut_FAT DEFAULT
    RESISTANCE 0.2700000000 ;
    LAYER M6 ;
        RECT -0.260 -0.260  0.260  0.260 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.260 -0.260  0.260  0.260 ;
END VIA67_1cut_FAT
                 
VIA VIA67_2cut_E DEFAULT
    RESISTANCE 0.1350000000 ;
    LAYER M6 ;
        RECT -0.200 -0.260  0.900  0.260 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT 0.520 -0.180  0.880  0.180 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.960  0.200 ;
END VIA67_2cut_E
VIA VIA67_2cut_W DEFAULT
    RESISTANCE 0.1350000000 ;
    LAYER M6 ;
        RECT -0.900 -0.260  0.200  0.260 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.880 -0.180  -0.520  0.180 ;
    LAYER M7 ;
        RECT -0.960 -0.200  0.260  0.200 ;
END VIA67_2cut_W
 
VIA VIA67_2cut_N DEFAULT
    RESISTANCE 0.1350000000 ;
    LAYER M6 ;
        RECT -0.200 -0.260  0.200  0.960 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.180 0.520  0.180  0.880 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.900 ;
END VIA67_2cut_N
 
VIA VIA67_2cut_S DEFAULT
    RESISTANCE 0.1350000000 ;
    LAYER M6 ;
        RECT -0.200 -0.960  0.200  0.260 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.180 -0.880  0.180  -0.520 ;
    LAYER M7 ;
        RECT -0.260 -0.900  0.260  0.200 ;
END VIA67_2cut_S
VIA VIA67_4cut DEFAULT
    RESISTANCE 0.0675000000 ;
    LAYER M6 ;
        RECT -0.650 -0.710  0.650  0.710 ;
    LAYER VIA6 ;
        RECT -0.630 -0.630  -0.270  -0.270 ;
        RECT -0.630 0.270  -0.270  0.630 ;
        RECT 0.270 0.270  0.630  0.630 ;
        RECT 0.270 -0.630  0.630  -0.270 ;
    LAYER M7 ;
        RECT -0.710 -0.650  0.710  0.650 ;
END VIA67_4cut
VIA VIA78_1cut DEFAULT
    RESISTANCE 0.2700000000 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.200  0.260 ;
END VIA78_1cut
VIA VIA78_1cut_H DEFAULT
    RESISTANCE 0.2700000000 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.260 -0.200  0.260  0.200 ;
END VIA78_1cut_H
                 
VIA VIA78_1cut_V DEFAULT
    RESISTANCE 0.2700000000 ;
    LAYER M7 ;
        RECT -0.200 -0.260  0.200  0.260 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.200  0.260 ;
END VIA78_1cut_V
VIA VIA78_1cut_FAT_C DEFAULT
    RESISTANCE 0.2700000000 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.200  0.260 ;
END VIA78_1cut_FAT_C
VIA VIA78_1cut_FAT_H DEFAULT
    RESISTANCE 0.2700000000 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.260 -0.200  0.260  0.200 ;
END VIA78_1cut_FAT_H
VIA VIA78_1cut_FAT_V DEFAULT
    RESISTANCE 0.2700000000 ;
    LAYER M7 ;
        RECT -0.200 -0.260  0.200  0.260 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.200  0.260 ;
END VIA78_1cut_FAT_V
VIA VIA78_1cut_FAT DEFAULT
    RESISTANCE 0.2700000000 ;
    LAYER M7 ;
        RECT -0.260 -0.260  0.260  0.260 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.260 -0.260  0.260  0.260 ;
END VIA78_1cut_FAT
VIA VIA78_1stack_E DEFAULT
    RESISTANCE 0.2700000000 ;
    LAYER M7 ;
        RECT -0.260 -0.200  1.155  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.200  0.260 ;
END VIA78_1stack_E
 
VIA VIA78_1stack_W DEFAULT
    RESISTANCE 0.2700000000 ;
    LAYER M7 ;
        RECT -1.155 -0.200  0.260  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.200  0.260 ;
END VIA78_1stack_W
                 
VIA VIA78_2cut_E DEFAULT
    RESISTANCE 0.1350000000 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.960  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT 0.520 -0.180  0.880  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.900  0.260 ;
END VIA78_2cut_E
VIA VIA78_2cut_W DEFAULT
    RESISTANCE 0.1350000000 ;
    LAYER M7 ;
        RECT -0.960 -0.200  0.260  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.880 -0.180  -0.520  0.180 ;
    LAYER M8 ;
        RECT -0.900 -0.260  0.200  0.260 ;
END VIA78_2cut_W
 
VIA VIA78_2cut_N DEFAULT
    RESISTANCE 0.1350000000 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.900 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.180 0.520  0.180  0.880 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.200  0.960 ;
END VIA78_2cut_N
 
VIA VIA78_2cut_S DEFAULT
    RESISTANCE 0.1350000000 ;
    LAYER M7 ;
        RECT -0.260 -0.900  0.260  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.180 -0.880  0.180  -0.520 ;
    LAYER M8 ;
        RECT -0.200 -0.960  0.200  0.260 ;
END VIA78_2cut_S
 
VIA VIA78_2stack_E DEFAULT
    RESISTANCE 0.1350000000 ;
    LAYER M7 ;
        RECT -0.260 -0.200  1.155  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT 0.520 -0.180  0.880  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.900  0.260 ;
END VIA78_2stack_E
VIA VIA78_2stack_W DEFAULT
    RESISTANCE 0.1350000000 ;
    LAYER M7 ;
        RECT -1.155 -0.200  0.260  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.880 -0.180  -0.520  0.180 ;
    LAYER M8 ;
        RECT -0.900 -0.260  0.200  0.260 ;
END VIA78_2stack_W
VIA VIA78_4cut DEFAULT
    RESISTANCE 0.0675000000 ;
    LAYER M7 ;
        RECT -0.710 -0.650  0.710  0.650 ;
    LAYER VIA7 ;
        RECT -0.630 -0.630  -0.270  -0.270 ;
        RECT -0.630 0.270  -0.270  0.630 ;
        RECT 0.270 0.270  0.630  0.630 ;
        RECT 0.270 -0.630  0.630  -0.270 ;
    LAYER M8 ;
        RECT -0.650 -0.710  0.650  0.710 ;
END VIA78_4cut
VIA VIA12_pin
    RESISTANCE 6.7000000000 ;
    LAYER M1 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER VIA1 ;
        RECT -0.035 -0.035  0.035  0.035 ;
    LAYER M2 ;
        RECT -0.035 -0.035  0.035  0.035 ;
END VIA12_pin
SITE core
    SIZE 0.140 BY 1.260 ;
    CLASS CORE ;
    SYMMETRY Y  ;
END core
SITE pad
    SIZE 0.140 BY 1.260 ;
    CLASS PAD ;
    SYMMETRY Y  ;
END pad
MACRO io
    SIZE 0.140 BY 1.260 ;
    CLASS PAD ;
    SYMMETRY X Y ;
END io
MACRO in01s01
    CLASS CORE ;
    FOREIGN in01s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.420 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.120 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.245 0.495 0.350 0.775 ;
        END
    END a
END in01s01
MACRO in01s02
    CLASS CORE ;
    FOREIGN in01s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.210 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.465 0.495 0.685 0.775 ;
        END
    END a
END in01s02
MACRO in01s03
    CLASS CORE ;
    FOREIGN in01s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.305 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.675 0.495 0.990 0.775 ;
        END
    END a
END in01s03
MACRO in01s04
    CLASS CORE ;
    FOREIGN in01s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.385 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.885 0.495 1.305 0.775 ;
        END
    END a
END in01s04
MACRO in01s06
    CLASS CORE ;
    FOREIGN in01s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.660 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.295 0.495 1.935 0.775 ;
        END
    END a
END in01s06
MACRO in01s08
    CLASS CORE ;
    FOREIGN in01s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.730 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.725 0.495 2.565 0.775 ;
        END
    END a
END in01s08
MACRO in01s10
    CLASS CORE ;
    FOREIGN in01s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 1.430 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.405 0.495 5.085 0.775 ;
        END
    END a
END in01s10
MACRO in01s20
    CLASS CORE ;
    FOREIGN in01s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 2.835 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.755 0.495 10.125 0.775 ;
        END
    END a
END in01s20
MACRO in01s40
    CLASS CORE ;
    FOREIGN in01s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 26.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 5.625 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.475 0.495 20.205 0.775 ;
        END
    END a
END in01s40
MACRO in01s80
    CLASS CORE ;
    FOREIGN in01s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 53.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 11.195 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 26.915 0.495 40.355 0.775 ;
        END
    END a
END in01s80
MACRO in01m01
    CLASS CORE ;
    FOREIGN in01m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.420 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.120 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.245 0.495 0.350 0.775 ;
        END
    END a
END in01m01
MACRO in01m02
    CLASS CORE ;
    FOREIGN in01m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.210 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.465 0.495 0.685 0.775 ;
        END
    END a
END in01m02
MACRO in01m03
    CLASS CORE ;
    FOREIGN in01m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.305 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.675 0.495 0.990 0.775 ;
        END
    END a
END in01m03
MACRO in01m04
    CLASS CORE ;
    FOREIGN in01m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.385 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.885 0.495 1.305 0.775 ;
        END
    END a
END in01m04
MACRO in01m06
    CLASS CORE ;
    FOREIGN in01m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.660 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.295 0.495 1.935 0.775 ;
        END
    END a
END in01m06
MACRO in01m08
    CLASS CORE ;
    FOREIGN in01m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.730 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.725 0.495 2.565 0.775 ;
        END
    END a
END in01m08
MACRO in01m10
    CLASS CORE ;
    FOREIGN in01m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 1.430 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.405 0.495 5.085 0.775 ;
        END
    END a
END in01m10
MACRO in01m20
    CLASS CORE ;
    FOREIGN in01m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 2.835 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.755 0.495 10.125 0.775 ;
        END
    END a
END in01m20
MACRO in01m40
    CLASS CORE ;
    FOREIGN in01m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 26.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 5.625 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.475 0.495 20.205 0.775 ;
        END
    END a
END in01m40
MACRO in01m80
    CLASS CORE ;
    FOREIGN in01m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 53.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 11.195 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 26.915 0.495 40.355 0.775 ;
        END
    END a
END in01m80
MACRO in01f01
    CLASS CORE ;
    FOREIGN in01f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.420 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.120 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.245 0.495 0.350 0.775 ;
        END
    END a
END in01f01
MACRO in01f02
    CLASS CORE ;
    FOREIGN in01f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.210 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.465 0.495 0.685 0.775 ;
        END
    END a
END in01f02
MACRO in01f03
    CLASS CORE ;
    FOREIGN in01f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.305 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.675 0.495 0.990 0.775 ;
        END
    END a
END in01f03
MACRO in01f04
    CLASS CORE ;
    FOREIGN in01f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.385 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.885 0.495 1.305 0.775 ;
        END
    END a
END in01f04
MACRO in01f06
    CLASS CORE ;
    FOREIGN in01f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.660 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.295 0.495 1.935 0.775 ;
        END
    END a
END in01f06
MACRO in01f08
    CLASS CORE ;
    FOREIGN in01f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.730 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.725 0.495 2.565 0.775 ;
        END
    END a
END in01f08
MACRO in01f10
    CLASS CORE ;
    FOREIGN in01f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 1.430 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.405 0.495 5.085 0.775 ;
        END
    END a
END in01f10
MACRO in01f20
    CLASS CORE ;
    FOREIGN in01f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 2.835 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.755 0.495 10.125 0.775 ;
        END
    END a
END in01f20
MACRO in01f40
    CLASS CORE ;
    FOREIGN in01f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 26.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 5.625 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.475 0.495 20.205 0.775 ;
        END
    END a
END in01f40
MACRO in01f80
    CLASS CORE ;
    FOREIGN in01f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 53.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 11.195 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 26.915 0.495 40.355 0.775 ;
        END
    END a
END in01f80
MACRO na02s01
    CLASS CORE ;
    FOREIGN na02s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.135 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.220 0.495 0.325 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.410 0.495 0.500 0.775 ;
        END
    END b
END na02s01
MACRO na02s02
    CLASS CORE ;
    FOREIGN na02s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.170 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.325 0.495 0.480 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.595 0.495 0.730 0.775 ;
        END
    END b
END na02s02
MACRO na02s03
    CLASS CORE ;
    FOREIGN na02s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.260 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.500 0.495 0.760 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.070 0.495 1.295 0.775 ;
        END
    END b
END na02s03
MACRO na02s04
    CLASS CORE ;
    FOREIGN na02s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.315 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.595 0.495 0.915 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.165 0.495 1.445 0.775 ;
        END
    END b
END na02s04
MACRO na02s06
    CLASS CORE ;
    FOREIGN na02s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.445 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.885 0.495 1.355 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.725 0.495 2.130 0.775 ;
        END
    END b
END na02s06
MACRO na02s08
    CLASS CORE ;
    FOREIGN na02s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.680 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.165 0.495 1.890 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.275 0.495 2.815 0.775 ;
        END
    END b
END na02s08
MACRO na02s10
    CLASS CORE ;
    FOREIGN na02s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 1.125 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.275 0.495 3.525 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.515 0.495 5.595 0.775 ;
        END
    END b
END na02s10
MACRO na02s20
    CLASS CORE ;
    FOREIGN na02s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 2.210 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.515 0.495 7.015 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.995 0.495 11.155 0.775 ;
        END
    END b
END na02s20
MACRO na02s40
    CLASS CORE ;
    FOREIGN na02s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 26.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 4.490 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.995 0.495 13.990 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 17.955 0.495 22.275 0.775 ;
        END
    END b
END na02s40
MACRO na02s80
    CLASS CORE ;
    FOREIGN na02s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 53.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 8.745 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 17.955 0.495 27.955 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 35.885 0.495 44.525 0.775 ;
        END
    END b
END na02s80
MACRO na02m01
    CLASS CORE ;
    FOREIGN na02m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.135 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.220 0.495 0.325 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.410 0.495 0.500 0.775 ;
        END
    END b
END na02m01
MACRO na02m02
    CLASS CORE ;
    FOREIGN na02m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.170 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.325 0.495 0.480 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.595 0.495 0.730 0.775 ;
        END
    END b
END na02m02
MACRO na02m03
    CLASS CORE ;
    FOREIGN na02m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.260 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.500 0.495 0.760 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.070 0.495 1.295 0.775 ;
        END
    END b
END na02m03
MACRO na02m04
    CLASS CORE ;
    FOREIGN na02m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.315 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.595 0.495 0.915 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.165 0.495 1.445 0.775 ;
        END
    END b
END na02m04
MACRO na02m06
    CLASS CORE ;
    FOREIGN na02m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.445 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.885 0.495 1.355 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.725 0.495 2.130 0.775 ;
        END
    END b
END na02m06
MACRO na02m08
    CLASS CORE ;
    FOREIGN na02m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.680 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.165 0.495 1.890 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.275 0.495 2.815 0.775 ;
        END
    END b
END na02m08
MACRO na02m10
    CLASS CORE ;
    FOREIGN na02m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 1.125 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.275 0.495 3.525 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.515 0.495 5.595 0.775 ;
        END
    END b
END na02m10
MACRO na02m20
    CLASS CORE ;
    FOREIGN na02m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 2.210 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.515 0.495 7.015 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.995 0.495 11.155 0.775 ;
        END
    END b
END na02m20
MACRO na02m40
    CLASS CORE ;
    FOREIGN na02m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 26.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 4.490 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.995 0.495 13.990 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 17.955 0.495 22.275 0.775 ;
        END
    END b
END na02m40
MACRO na02m80
    CLASS CORE ;
    FOREIGN na02m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 53.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 8.745 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 17.955 0.495 27.955 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 35.885 0.495 44.525 0.775 ;
        END
    END b
END na02m80
MACRO na02f01
    CLASS CORE ;
    FOREIGN na02f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.135 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.220 0.495 0.325 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.410 0.495 0.500 0.775 ;
        END
    END b
END na02f01
MACRO na02f02
    CLASS CORE ;
    FOREIGN na02f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.170 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.325 0.495 0.480 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.595 0.495 0.730 0.775 ;
        END
    END b
END na02f02
MACRO na02f03
    CLASS CORE ;
    FOREIGN na02f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.260 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.500 0.495 0.760 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.070 0.495 1.295 0.775 ;
        END
    END b
END na02f03
MACRO na02f04
    CLASS CORE ;
    FOREIGN na02f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.315 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.595 0.495 0.915 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.165 0.495 1.445 0.775 ;
        END
    END b
END na02f04
MACRO na02f06
    CLASS CORE ;
    FOREIGN na02f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.445 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.885 0.495 1.355 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.725 0.495 2.130 0.775 ;
        END
    END b
END na02f06
MACRO na02f08
    CLASS CORE ;
    FOREIGN na02f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.680 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.165 0.495 1.890 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.275 0.495 2.815 0.775 ;
        END
    END b
END na02f08
MACRO na02f10
    CLASS CORE ;
    FOREIGN na02f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 1.125 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.275 0.495 3.525 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.515 0.495 5.595 0.775 ;
        END
    END b
END na02f10
MACRO na02f20
    CLASS CORE ;
    FOREIGN na02f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 2.210 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.515 0.495 7.015 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.995 0.495 11.155 0.775 ;
        END
    END b
END na02f20
MACRO na02f40
    CLASS CORE ;
    FOREIGN na02f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 26.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 4.490 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.995 0.495 13.990 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 17.955 0.495 22.275 0.775 ;
        END
    END b
END na02f40
MACRO na02f80
    CLASS CORE ;
    FOREIGN na02f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 53.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 8.745 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 17.955 0.495 27.955 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 35.885 0.495 44.525 0.775 ;
        END
    END b
END na02f80
MACRO na03s01
    CLASS CORE ;
    FOREIGN na03s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 0.205 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.245 0.495 0.350 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.465 0.570 0.545 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.675 0.410 0.880 0.850 ;
        END
    END c
END na03s01
MACRO na03s02
    CLASS CORE ;
    FOREIGN na03s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 0.285 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.350 0.495 0.515 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.675 0.570 0.785 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.980 0.410 1.135 0.850 ;
        END
    END c
END na03s02
MACRO na03s03
    CLASS CORE ;
    FOREIGN na03s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 0.365 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.465 0.495 0.675 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.885 0.570 1.030 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.295 0.410 1.500 0.850 ;
        END
    END c
END na03s03
MACRO na03s04
    CLASS CORE ;
    FOREIGN na03s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 0.525 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.675 0.495 0.995 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.295 0.570 1.510 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.935 0.410 2.245 0.850 ;
        END
    END c
END na03s04
MACRO na03s06
    CLASS CORE ;
    FOREIGN na03s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 0.685 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.885 0.495 1.300 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.725 0.570 2.015 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.565 0.410 2.985 0.850 ;
        END
    END c
END na03s06
MACRO na03s08
    CLASS CORE ;
    FOREIGN na03s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 0.920 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.190 0.495 1.760 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.355 0.570 2.750 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.500 0.410 4.075 0.850 ;
        END
    END c
END na03s08
MACRO na03s10
    CLASS CORE ;
    FOREIGN na03s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 1.800 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.355 0.495 3.500 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.665 0.570 5.465 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.965 0.410 8.105 0.850 ;
        END
    END c
END na03s10
MACRO na03s20
    CLASS CORE ;
    FOREIGN na03s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 3.590 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.550 0.495 6.890 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 9.065 0.570 10.615 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.580 0.410 15.890 0.850 ;
        END
    END c
END na03s20
MACRO na03s40
    CLASS CORE ;
    FOREIGN na03s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 36.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 6.940 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 9.065 0.495 13.540 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 18.095 0.570 21.190 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 27.125 0.410 31.545 0.850 ;
        END
    END c
END na03s40
MACRO na03s80
    CLASS CORE ;
    FOREIGN na03s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 71.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 13.775 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 17.990 0.495 26.990 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 35.955 0.570 42.110 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 53.900 0.410 62.695 0.850 ;
        END
    END c
END na03s80
MACRO na03m01
    CLASS CORE ;
    FOREIGN na03m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 0.205 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.245 0.495 0.350 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.465 0.570 0.545 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.675 0.410 0.880 0.850 ;
        END
    END c
END na03m01
MACRO na03m02
    CLASS CORE ;
    FOREIGN na03m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 0.285 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.350 0.495 0.515 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.675 0.570 0.785 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.980 0.410 1.135 0.850 ;
        END
    END c
END na03m02
MACRO na03m03
    CLASS CORE ;
    FOREIGN na03m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 0.365 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.465 0.495 0.675 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.885 0.570 1.030 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.295 0.410 1.500 0.850 ;
        END
    END c
END na03m03
MACRO na03m04
    CLASS CORE ;
    FOREIGN na03m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 0.525 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.675 0.495 0.995 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.295 0.570 1.510 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.935 0.410 2.245 0.850 ;
        END
    END c
END na03m04
MACRO na03m06
    CLASS CORE ;
    FOREIGN na03m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 0.685 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.885 0.495 1.300 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.725 0.570 2.015 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.565 0.410 2.985 0.850 ;
        END
    END c
END na03m06
MACRO na03m08
    CLASS CORE ;
    FOREIGN na03m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 0.920 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.190 0.495 1.760 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.355 0.570 2.750 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.500 0.410 4.075 0.850 ;
        END
    END c
END na03m08
MACRO na03m10
    CLASS CORE ;
    FOREIGN na03m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 1.800 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.355 0.495 3.500 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.665 0.570 5.465 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.965 0.410 8.105 0.850 ;
        END
    END c
END na03m10
MACRO na03m20
    CLASS CORE ;
    FOREIGN na03m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 3.590 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.550 0.495 6.890 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 9.065 0.570 10.615 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.580 0.410 15.890 0.850 ;
        END
    END c
END na03m20
MACRO na03m40
    CLASS CORE ;
    FOREIGN na03m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 36.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 6.940 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 9.065 0.495 13.540 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 18.095 0.570 21.190 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 27.125 0.410 31.545 0.850 ;
        END
    END c
END na03m40
MACRO na03m80
    CLASS CORE ;
    FOREIGN na03m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 71.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 13.775 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 17.990 0.495 26.990 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 35.955 0.570 42.110 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 53.900 0.410 62.695 0.850 ;
        END
    END c
END na03m80
MACRO na03f01
    CLASS CORE ;
    FOREIGN na03f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 0.205 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.245 0.495 0.350 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.465 0.570 0.545 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.675 0.410 0.880 0.850 ;
        END
    END c
END na03f01
MACRO na03f02
    CLASS CORE ;
    FOREIGN na03f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 0.285 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.350 0.495 0.515 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.675 0.570 0.785 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.980 0.410 1.135 0.850 ;
        END
    END c
END na03f02
MACRO na03f03
    CLASS CORE ;
    FOREIGN na03f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 0.365 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.465 0.495 0.675 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.885 0.570 1.030 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.295 0.410 1.500 0.850 ;
        END
    END c
END na03f03
MACRO na03f04
    CLASS CORE ;
    FOREIGN na03f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 0.525 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.675 0.495 0.995 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.295 0.570 1.510 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.935 0.410 2.245 0.850 ;
        END
    END c
END na03f04
MACRO na03f06
    CLASS CORE ;
    FOREIGN na03f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 0.685 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.885 0.495 1.300 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.725 0.570 2.015 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.565 0.410 2.985 0.850 ;
        END
    END c
END na03f06
MACRO na03f08
    CLASS CORE ;
    FOREIGN na03f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 0.920 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.190 0.495 1.760 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.355 0.570 2.750 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.500 0.410 4.075 0.850 ;
        END
    END c
END na03f08
MACRO na03f10
    CLASS CORE ;
    FOREIGN na03f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 1.800 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.355 0.495 3.500 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.665 0.570 5.465 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.965 0.410 8.105 0.850 ;
        END
    END c
END na03f10
MACRO na03f20
    CLASS CORE ;
    FOREIGN na03f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 3.590 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.550 0.495 6.890 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 9.065 0.570 10.615 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.580 0.410 15.890 0.850 ;
        END
    END c
END na03f20
MACRO na03f40
    CLASS CORE ;
    FOREIGN na03f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 36.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 6.940 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 9.065 0.495 13.540 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 18.095 0.570 21.190 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 27.125 0.410 31.545 0.850 ;
        END
    END c
END na03f40
MACRO na03f80
    CLASS CORE ;
    FOREIGN na03f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 71.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.290 13.775 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 17.990 0.495 26.990 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 35.955 0.570 42.110 0.790 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 53.900 0.410 62.695 0.850 ;
        END
    END c
END na03f80
MACRO na04s01
    CLASS CORE ;
    FOREIGN na04s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 0.195 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.230 0.495 0.340 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.435 0.475 0.515 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.625 0.495 0.730 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.820 0.475 0.890 0.795 ;
        END
    END d
END na04s01
MACRO na04s02
    CLASS CORE ;
    FOREIGN na04s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.470 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 0.260 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.330 0.495 0.505 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.625 0.475 0.730 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.925 0.495 1.080 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.210 0.475 1.315 0.795 ;
        END
    END d
END na04s02
MACRO na04s03
    CLASS CORE ;
    FOREIGN na04s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 0.340 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.435 0.495 0.760 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.820 0.475 0.960 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.210 0.495 1.420 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.605 0.475 1.755 0.795 ;
        END
    END d
END na04s03
MACRO na04s04
    CLASS CORE ;
    FOREIGN na04s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.450 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 0.415 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.535 0.495 0.815 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.015 0.475 1.190 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.495 1.765 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.475 2.180 0.795 ;
        END
    END d
END na04s04
MACRO na04s06
    CLASS CORE ;
    FOREIGN na04s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 0.640 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.820 0.495 1.275 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.605 0.475 1.895 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.395 0.495 2.810 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.170 0.475 3.450 0.795 ;
        END
    END d
END na04s06
MACRO na04s08
    CLASS CORE ;
    FOREIGN na04s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 0.795 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.015 0.495 1.570 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.475 2.355 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.985 0.495 3.505 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.475 4.325 0.795 ;
        END
    END d
END na04s08
MACRO na04s10
    CLASS CORE ;
    FOREIGN na04s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 1.550 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.495 3.120 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.475 4.675 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.925 0.495 6.975 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.475 8.595 0.795 ;
        END
    END d
END na04s10
MACRO na04s20
    CLASS CORE ;
    FOREIGN na04s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 3.065 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.495 6.205 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.475 9.295 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 11.795 0.495 13.885 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.475 17.115 0.795 ;
        END
    END d
END na04s20
MACRO na04s40
    CLASS CORE ;
    FOREIGN na04s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 39.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 6.105 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.495 12.345 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.475 18.525 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 23.555 0.495 27.720 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 31.395 0.475 34.205 0.795 ;
        END
    END d
END na04s40
MACRO na04s80
    CLASS CORE ;
    FOREIGN na04s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 78.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 12.165 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.495 24.635 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 31.395 0.475 36.995 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 47.085 0.495 55.410 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 62.765 0.475 68.365 0.795 ;
        END
    END d
END na04s80
MACRO na04m01
    CLASS CORE ;
    FOREIGN na04m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 0.195 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.230 0.495 0.340 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.435 0.475 0.515 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.625 0.495 0.730 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.820 0.475 0.890 0.795 ;
        END
    END d
END na04m01
MACRO na04m02
    CLASS CORE ;
    FOREIGN na04m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.470 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 0.260 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.330 0.495 0.505 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.625 0.475 0.730 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.925 0.495 1.080 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.210 0.475 1.315 0.795 ;
        END
    END d
END na04m02
MACRO na04m03
    CLASS CORE ;
    FOREIGN na04m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 0.340 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.435 0.495 0.760 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.820 0.475 0.960 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.210 0.495 1.420 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.605 0.475 1.755 0.795 ;
        END
    END d
END na04m03
MACRO na04m04
    CLASS CORE ;
    FOREIGN na04m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.450 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 0.415 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.535 0.495 0.815 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.015 0.475 1.190 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.495 1.765 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.475 2.180 0.795 ;
        END
    END d
END na04m04
MACRO na04m06
    CLASS CORE ;
    FOREIGN na04m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 0.640 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.820 0.495 1.275 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.605 0.475 1.895 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.395 0.495 2.810 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.170 0.475 3.450 0.795 ;
        END
    END d
END na04m06
MACRO na04m08
    CLASS CORE ;
    FOREIGN na04m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 0.795 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.015 0.495 1.570 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.475 2.355 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.985 0.495 3.505 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.475 4.325 0.795 ;
        END
    END d
END na04m08
MACRO na04m10
    CLASS CORE ;
    FOREIGN na04m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 1.550 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.495 3.120 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.475 4.675 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.925 0.495 6.975 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.475 8.595 0.795 ;
        END
    END d
END na04m10
MACRO na04m20
    CLASS CORE ;
    FOREIGN na04m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 3.065 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.495 6.205 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.475 9.295 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 11.795 0.495 13.885 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.475 17.115 0.795 ;
        END
    END d
END na04m20
MACRO na04m40
    CLASS CORE ;
    FOREIGN na04m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 39.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 6.105 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.495 12.345 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.475 18.525 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 23.555 0.495 27.720 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 31.395 0.475 34.205 0.795 ;
        END
    END d
END na04m40
MACRO na04m80
    CLASS CORE ;
    FOREIGN na04m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 78.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 12.165 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.495 24.635 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 31.395 0.475 36.995 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 47.085 0.495 55.410 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 62.765 0.475 68.365 0.795 ;
        END
    END d
END na04m80
MACRO na04f01
    CLASS CORE ;
    FOREIGN na04f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 0.195 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.230 0.495 0.340 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.435 0.475 0.515 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.625 0.495 0.730 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.820 0.475 0.890 0.795 ;
        END
    END d
END na04f01
MACRO na04f02
    CLASS CORE ;
    FOREIGN na04f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.470 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 0.260 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.330 0.495 0.505 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.625 0.475 0.730 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.925 0.495 1.080 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.210 0.475 1.315 0.795 ;
        END
    END d
END na04f02
MACRO na04f03
    CLASS CORE ;
    FOREIGN na04f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 0.340 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.435 0.495 0.760 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.820 0.475 0.960 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.210 0.495 1.420 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.605 0.475 1.755 0.795 ;
        END
    END d
END na04f03
MACRO na04f04
    CLASS CORE ;
    FOREIGN na04f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.450 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 0.415 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.535 0.495 0.815 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.015 0.475 1.190 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.495 1.765 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.475 2.180 0.795 ;
        END
    END d
END na04f04
MACRO na04f06
    CLASS CORE ;
    FOREIGN na04f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 0.640 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.820 0.495 1.275 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.605 0.475 1.895 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.395 0.495 2.810 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.170 0.475 3.450 0.795 ;
        END
    END d
END na04f06
MACRO na04f08
    CLASS CORE ;
    FOREIGN na04f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 0.795 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.015 0.495 1.570 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.475 2.355 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.985 0.495 3.505 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.475 4.325 0.795 ;
        END
    END d
END na04f08
MACRO na04f10
    CLASS CORE ;
    FOREIGN na04f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 1.550 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.495 3.120 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.475 4.675 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.925 0.495 6.975 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.475 8.595 0.795 ;
        END
    END d
END na04f10
MACRO na04f20
    CLASS CORE ;
    FOREIGN na04f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 3.065 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.495 6.205 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.475 9.295 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 11.795 0.495 13.885 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.475 17.115 0.795 ;
        END
    END d
END na04f20
MACRO na04f40
    CLASS CORE ;
    FOREIGN na04f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 39.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 6.105 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.495 12.345 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.475 18.525 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 23.555 0.495 27.720 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 31.395 0.475 34.205 0.795 ;
        END
    END d
END na04f40
MACRO na04f80
    CLASS CORE ;
    FOREIGN na04f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 78.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.210 12.165 1.050 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.495 24.635 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 31.395 0.475 36.995 0.795 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 47.085 0.495 55.410 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 62.765 0.475 68.365 0.795 ;
        END
    END d
END na04f80
MACRO no02s01
    CLASS CORE ;
    FOREIGN no02s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.135 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.220 0.590 0.330 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.410 0.495 0.500 0.775 ;
        END
    END b
END no02s01
MACRO no02s02
    CLASS CORE ;
    FOREIGN no02s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.170 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.325 0.590 0.495 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.595 0.495 0.730 0.775 ;
        END
    END b
END no02s02
MACRO no02s03
    CLASS CORE ;
    FOREIGN no02s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.260 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.500 0.590 0.770 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.070 0.495 1.295 0.775 ;
        END
    END b
END no02s03
MACRO no02s04
    CLASS CORE ;
    FOREIGN no02s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.315 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.595 0.590 0.920 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.165 0.495 1.445 0.775 ;
        END
    END b
END no02s04
MACRO no02s06
    CLASS CORE ;
    FOREIGN no02s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.445 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.885 0.590 1.370 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.725 0.495 2.130 0.775 ;
        END
    END b
END no02s06
MACRO no02s08
    CLASS CORE ;
    FOREIGN no02s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.680 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.165 0.590 1.810 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.275 0.495 2.815 0.775 ;
        END
    END b
END no02s08
MACRO no02s10
    CLASS CORE ;
    FOREIGN no02s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 1.125 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.275 0.590 3.570 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.515 0.495 5.595 0.775 ;
        END
    END b
END no02s10
MACRO no02s20
    CLASS CORE ;
    FOREIGN no02s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 2.210 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.515 0.590 7.105 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.995 0.495 11.155 0.775 ;
        END
    END b
END no02s20
MACRO no02s40
    CLASS CORE ;
    FOREIGN no02s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 26.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 4.490 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.995 0.590 14.175 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 17.955 0.495 22.275 0.775 ;
        END
    END b
END no02s40
MACRO no02s80
    CLASS CORE ;
    FOREIGN no02s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 53.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 8.745 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 17.955 0.590 28.315 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 35.885 0.495 44.525 0.775 ;
        END
    END b
END no02s80
MACRO no02m01
    CLASS CORE ;
    FOREIGN no02m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.135 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.220 0.590 0.330 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.410 0.495 0.500 0.775 ;
        END
    END b
END no02m01
MACRO no02m02
    CLASS CORE ;
    FOREIGN no02m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.170 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.325 0.590 0.495 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.595 0.495 0.730 0.775 ;
        END
    END b
END no02m02
MACRO no02m03
    CLASS CORE ;
    FOREIGN no02m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.260 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.500 0.590 0.770 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.070 0.495 1.295 0.775 ;
        END
    END b
END no02m03
MACRO no02m04
    CLASS CORE ;
    FOREIGN no02m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.315 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.595 0.590 0.920 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.165 0.495 1.445 0.775 ;
        END
    END b
END no02m04
MACRO no02m06
    CLASS CORE ;
    FOREIGN no02m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.445 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.885 0.590 1.370 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.725 0.495 2.130 0.775 ;
        END
    END b
END no02m06
MACRO no02m08
    CLASS CORE ;
    FOREIGN no02m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.680 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.165 0.590 1.810 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.275 0.495 2.815 0.775 ;
        END
    END b
END no02m08
MACRO no02m10
    CLASS CORE ;
    FOREIGN no02m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 1.125 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.275 0.590 3.570 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.515 0.495 5.595 0.775 ;
        END
    END b
END no02m10
MACRO no02m20
    CLASS CORE ;
    FOREIGN no02m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 2.210 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.515 0.590 7.105 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.995 0.495 11.155 0.775 ;
        END
    END b
END no02m20
MACRO no02m40
    CLASS CORE ;
    FOREIGN no02m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 26.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 4.490 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.995 0.590 14.175 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 17.955 0.495 22.275 0.775 ;
        END
    END b
END no02m40
MACRO no02m80
    CLASS CORE ;
    FOREIGN no02m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 53.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 8.745 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 17.955 0.590 28.315 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 35.885 0.495 44.525 0.775 ;
        END
    END b
END no02m80
MACRO no02f01
    CLASS CORE ;
    FOREIGN no02f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.135 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.220 0.590 0.330 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.410 0.495 0.500 0.775 ;
        END
    END b
END no02f01
MACRO no02f02
    CLASS CORE ;
    FOREIGN no02f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.170 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.325 0.590 0.495 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.595 0.495 0.730 0.775 ;
        END
    END b
END no02f02
MACRO no02f03
    CLASS CORE ;
    FOREIGN no02f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.260 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.500 0.590 0.770 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.070 0.495 1.295 0.775 ;
        END
    END b
END no02f03
MACRO no02f04
    CLASS CORE ;
    FOREIGN no02f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.315 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.595 0.590 0.920 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.165 0.495 1.445 0.775 ;
        END
    END b
END no02f04
MACRO no02f06
    CLASS CORE ;
    FOREIGN no02f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.445 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.885 0.590 1.370 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.725 0.495 2.130 0.775 ;
        END
    END b
END no02f06
MACRO no02f08
    CLASS CORE ;
    FOREIGN no02f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 0.680 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.165 0.590 1.810 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.275 0.495 2.815 0.775 ;
        END
    END b
END no02f08
MACRO no02f10
    CLASS CORE ;
    FOREIGN no02f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 1.125 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.275 0.590 3.570 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.515 0.495 5.595 0.775 ;
        END
    END b
END no02f10
MACRO no02f20
    CLASS CORE ;
    FOREIGN no02f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 2.210 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.515 0.590 7.105 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.995 0.495 11.155 0.775 ;
        END
    END b
END no02f20
MACRO no02f40
    CLASS CORE ;
    FOREIGN no02f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 26.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 4.490 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.995 0.590 14.175 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 17.955 0.495 22.275 0.775 ;
        END
    END b
END no02f40
MACRO no02f80
    CLASS CORE ;
    FOREIGN no02f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 53.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.215 8.745 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 17.955 0.590 28.315 0.770 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 35.885 0.495 44.525 0.775 ;
        END
    END b
END no02f80
MACRO no03s01
    CLASS CORE ;
    FOREIGN no03s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 0.310 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.350 0.565 0.560 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.675 0.590 0.905 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.980 0.405 1.225 0.865 ;
        END
    END c
END no03s01
MACRO no03s02
    CLASS CORE ;
    FOREIGN no03s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.890 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 0.450 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.510 0.565 0.825 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.980 0.590 1.310 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.450 0.405 1.825 0.865 ;
        END
    END c
END no03s02
MACRO no03s03
    CLASS CORE ;
    FOREIGN no03s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 0.595 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.675 0.565 1.095 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.295 0.590 1.745 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.935 0.405 2.425 0.865 ;
        END
    END c
END no03s03
MACRO no03s04
    CLASS CORE ;
    FOREIGN no03s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 0.860 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.980 0.565 1.610 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.935 0.590 2.6100 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.870 0.405 3.600 0.865 ;
        END
    END c
END no03s04
MACRO no03s06
    CLASS CORE ;
    FOREIGN no03s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 1.140 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.295 0.565 2.135 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.565 0.590 3.450 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.815 0.405 4.790 0.865 ;
        END
    END c
END no03s06
MACRO no03s08
    CLASS CORE ;
    FOREIGN no03s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 1.550 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.775 0.565 2.930 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.500 0.590 4.725 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.235 0.405 6.585 0.865 ;
        END
    END c
END no03s08
MACRO no03s10
    CLASS CORE ;
    FOREIGN no03s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 3.075 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.500 0.565 5.810 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.965 0.590 9.405 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 10.430 0.405 13.110 0.865 ;
        END
    END c
END no03s10
MACRO no03s20
    CLASS CORE ;
    FOREIGN no03s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 27.090 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 5.960 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.810 0.565 11.325 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.580 0.590 18.335 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 20.355 0.405 25.605 0.865 ;
        END
    END c
END no03s20
MACRO no03s40
    CLASS CORE ;
    FOREIGN no03s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 54.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 11.990 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.580 0.565 22.610 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 27.125 0.590 36.630 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 40.670 0.405 51.155 0.865 ;
        END
    END c
END no03s40
MACRO no03s80
    CLASS CORE ;
    FOREIGN no03s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 107.730 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 23.605 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 27.070 0.565 45.025 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 53.900 0.590 72.800 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 80.830 0.405 101.685 0.865 ;
        END
    END c
END no03s80
MACRO no03m01
    CLASS CORE ;
    FOREIGN no03m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 0.310 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.350 0.565 0.560 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.675 0.590 0.905 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.980 0.405 1.225 0.865 ;
        END
    END c
END no03m01
MACRO no03m02
    CLASS CORE ;
    FOREIGN no03m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.890 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 0.450 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.510 0.565 0.825 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.980 0.590 1.310 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.450 0.405 1.825 0.865 ;
        END
    END c
END no03m02
MACRO no03m03
    CLASS CORE ;
    FOREIGN no03m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 0.595 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.675 0.565 1.095 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.295 0.590 1.745 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.935 0.405 2.425 0.865 ;
        END
    END c
END no03m03
MACRO no03m04
    CLASS CORE ;
    FOREIGN no03m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 0.860 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.980 0.565 1.610 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.935 0.590 2.6100 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.870 0.405 3.600 0.865 ;
        END
    END c
END no03m04
MACRO no03m06
    CLASS CORE ;
    FOREIGN no03m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 1.140 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.295 0.565 2.135 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.565 0.590 3.450 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.815 0.405 4.790 0.865 ;
        END
    END c
END no03m06
MACRO no03m08
    CLASS CORE ;
    FOREIGN no03m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 1.550 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.775 0.565 2.930 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.500 0.590 4.725 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.235 0.405 6.585 0.865 ;
        END
    END c
END no03m08
MACRO no03m10
    CLASS CORE ;
    FOREIGN no03m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 3.075 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.500 0.565 5.810 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.965 0.590 9.405 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 10.430 0.405 13.110 0.865 ;
        END
    END c
END no03m10
MACRO no03m20
    CLASS CORE ;
    FOREIGN no03m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 27.090 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 5.960 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.810 0.565 11.325 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.580 0.590 18.335 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 20.355 0.405 25.605 0.865 ;
        END
    END c
END no03m20
MACRO no03m40
    CLASS CORE ;
    FOREIGN no03m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 54.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 11.990 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.580 0.565 22.610 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 27.125 0.590 36.630 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 40.670 0.405 51.155 0.865 ;
        END
    END c
END no03m40
MACRO no03m80
    CLASS CORE ;
    FOREIGN no03m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 107.730 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 23.605 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 27.070 0.565 45.025 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 53.900 0.590 72.800 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 80.830 0.405 101.685 0.865 ;
        END
    END c
END no03m80
MACRO no03f01
    CLASS CORE ;
    FOREIGN no03f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 0.310 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.350 0.565 0.560 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.675 0.590 0.905 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.980 0.405 1.225 0.865 ;
        END
    END c
END no03f01
MACRO no03f02
    CLASS CORE ;
    FOREIGN no03f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.890 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 0.450 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.510 0.565 0.825 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.980 0.590 1.310 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.450 0.405 1.825 0.865 ;
        END
    END c
END no03f02
MACRO no03f03
    CLASS CORE ;
    FOREIGN no03f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 0.595 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.675 0.565 1.095 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.295 0.590 1.745 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.935 0.405 2.425 0.865 ;
        END
    END c
END no03f03
MACRO no03f04
    CLASS CORE ;
    FOREIGN no03f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 0.860 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.980 0.565 1.610 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.935 0.590 2.6100 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.870 0.405 3.600 0.865 ;
        END
    END c
END no03f04
MACRO no03f06
    CLASS CORE ;
    FOREIGN no03f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 1.140 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.295 0.565 2.135 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.565 0.590 3.450 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.815 0.405 4.790 0.865 ;
        END
    END c
END no03f06
MACRO no03f08
    CLASS CORE ;
    FOREIGN no03f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.930 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 1.550 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.775 0.565 2.930 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.500 0.590 4.725 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.235 0.405 6.585 0.865 ;
        END
    END c
END no03f08
MACRO no03f10
    CLASS CORE ;
    FOREIGN no03f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.860 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 3.075 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.500 0.565 5.810 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.965 0.590 9.405 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 10.430 0.405 13.110 0.865 ;
        END
    END c
END no03f10
MACRO no03f20
    CLASS CORE ;
    FOREIGN no03f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 27.090 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 5.960 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.810 0.565 11.325 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.580 0.590 18.335 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 20.355 0.405 25.605 0.865 ;
        END
    END c
END no03f20
MACRO no03f40
    CLASS CORE ;
    FOREIGN no03f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 54.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 11.990 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.580 0.565 22.610 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 27.125 0.590 36.630 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 40.670 0.405 51.155 0.865 ;
        END
    END c
END no03f40
MACRO no03f80
    CLASS CORE ;
    FOREIGN no03f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 107.730 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.2100 23.605 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 27.070 0.565 45.025 0.695 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 53.900 0.590 72.800 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 80.830 0.405 101.685 0.865 ;
        END
    END c
END no03f80
MACRO no04s01
    CLASS CORE ;
    FOREIGN no04s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 0.330 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.370 0.495 0.455 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.715 0.495 0.8100 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.490 1.160 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.480 0.590 1.565 0.770 ;
        END
    END d
END no04s01
MACRO no04s02
    CLASS CORE ;
    FOREIGN no04s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 0.485 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.540 0.495 0.675 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.495 1.170 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.490 1.730 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.590 2.175 0.770 ;
        END
    END d
END no04s02
MACRO no04s03
    CLASS CORE ;
    FOREIGN no04s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 0.625 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.715 0.495 0.880 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.480 0.495 1.655 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.490 2.295 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.725 0.590 2.890 0.770 ;
        END
    END d
END no04s03
MACRO no04s04
    CLASS CORE ;
    FOREIGN no04s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 0.770 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.885 0.495 1.095 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.725 0.495 1.935 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.565 0.490 2.960 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.405 0.590 3.615 0.770 ;
        END
    END d
END no04s04
MACRO no04s06
    CLASS CORE ;
    FOREIGN no04s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 1.215 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.480 0.495 1.815 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.725 0.495 3.160 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.490 4.545 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.410 0.590 5.745 0.770 ;
        END
    END d
END no04s06
MACRO no04s08
    CLASS CORE ;
    FOREIGN no04s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 1.510 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.725 0.495 2.140 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.405 0.495 3.820 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.085 0.490 5.670 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.755 0.590 7.170 0.770 ;
        END
    END d
END no04s08
MACRO no04s10
    CLASS CORE ;
    FOREIGN no04s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 2.985 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.405 0.495 4.240 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.755 0.495 7.690 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 10.125 0.490 11.3100 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.475 0.590 14.310 0.770 ;
        END
    END d
END no04s10
MACRO no04s20
    CLASS CORE ;
    FOREIGN no04s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 33.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 5.930 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.755 0.495 8.425 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.475 0.495 15.145 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 20.205 0.490 22.550 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 26.915 0.590 28.585 0.770 ;
        END
    END d
END no04s20
MACRO no04s40
    CLASS CORE ;
    FOREIGN no04s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 67.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 11.835 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.475 0.495 16.810 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 26.915 0.495 30.250 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 40.355 0.490 45.055 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 53.805 0.590 57.140 0.770 ;
        END
    END d
END no04s40
MACRO no04s80
    CLASS CORE ;
    FOREIGN no04s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 134.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 23.625 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 26.915 0.495 33.690 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 53.805 0.495 60.580 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 80.675 0.490 90.065 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 107.565 0.590 114.240 0.770 ;
        END
    END d
END no04s80
MACRO no04m01
    CLASS CORE ;
    FOREIGN no04m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 0.330 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.370 0.495 0.455 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.715 0.495 0.8100 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.490 1.160 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.480 0.590 1.565 0.770 ;
        END
    END d
END no04m01
MACRO no04m02
    CLASS CORE ;
    FOREIGN no04m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 0.485 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.540 0.495 0.675 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.495 1.170 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.490 1.730 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.590 2.175 0.770 ;
        END
    END d
END no04m02
MACRO no04m03
    CLASS CORE ;
    FOREIGN no04m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 0.625 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.715 0.495 0.880 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.480 0.495 1.655 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.490 2.295 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.725 0.590 2.890 0.770 ;
        END
    END d
END no04m03
MACRO no04m04
    CLASS CORE ;
    FOREIGN no04m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 0.770 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.885 0.495 1.095 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.725 0.495 1.935 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.565 0.490 2.960 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.405 0.590 3.615 0.770 ;
        END
    END d
END no04m04
MACRO no04m06
    CLASS CORE ;
    FOREIGN no04m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 1.215 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.480 0.495 1.815 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.725 0.495 3.160 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.490 4.545 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.410 0.590 5.745 0.770 ;
        END
    END d
END no04m06
MACRO no04m08
    CLASS CORE ;
    FOREIGN no04m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 1.510 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.725 0.495 2.140 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.405 0.495 3.820 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.085 0.490 5.670 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.755 0.590 7.170 0.770 ;
        END
    END d
END no04m08
MACRO no04m10
    CLASS CORE ;
    FOREIGN no04m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 2.985 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.405 0.495 4.240 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.755 0.495 7.690 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 10.125 0.490 11.3100 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.475 0.590 14.310 0.770 ;
        END
    END d
END no04m10
MACRO no04m20
    CLASS CORE ;
    FOREIGN no04m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 33.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 5.930 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.755 0.495 8.425 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.475 0.495 15.145 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 20.205 0.490 22.550 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 26.915 0.590 28.585 0.770 ;
        END
    END d
END no04m20
MACRO no04m40
    CLASS CORE ;
    FOREIGN no04m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 67.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 11.835 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.475 0.495 16.810 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 26.915 0.495 30.250 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 40.355 0.490 45.055 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 53.805 0.590 57.140 0.770 ;
        END
    END d
END no04m40
MACRO no04m80
    CLASS CORE ;
    FOREIGN no04m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 134.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 23.625 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 26.915 0.495 33.690 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 53.805 0.495 60.580 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 80.675 0.490 90.065 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 107.565 0.590 114.240 0.770 ;
        END
    END d
END no04m80
MACRO no04f01
    CLASS CORE ;
    FOREIGN no04f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 0.330 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.370 0.495 0.455 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.715 0.495 0.8100 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.490 1.160 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.480 0.590 1.565 0.770 ;
        END
    END d
END no04f01
MACRO no04f02
    CLASS CORE ;
    FOREIGN no04f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 0.485 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.540 0.495 0.675 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.495 1.170 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.490 1.730 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.590 2.175 0.770 ;
        END
    END d
END no04f02
MACRO no04f03
    CLASS CORE ;
    FOREIGN no04f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 0.625 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.715 0.495 0.880 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.480 0.495 1.655 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.490 2.295 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.725 0.590 2.890 0.770 ;
        END
    END d
END no04f03
MACRO no04f04
    CLASS CORE ;
    FOREIGN no04f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 0.770 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.885 0.495 1.095 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.725 0.495 1.935 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.565 0.490 2.960 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.405 0.590 3.615 0.770 ;
        END
    END d
END no04f04
MACRO no04f06
    CLASS CORE ;
    FOREIGN no04f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 1.215 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.480 0.495 1.815 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.725 0.495 3.160 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.490 4.545 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.410 0.590 5.745 0.770 ;
        END
    END d
END no04f06
MACRO no04f08
    CLASS CORE ;
    FOREIGN no04f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 1.510 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.725 0.495 2.140 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.405 0.495 3.820 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.085 0.490 5.670 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.755 0.590 7.170 0.770 ;
        END
    END d
END no04f08
MACRO no04f10
    CLASS CORE ;
    FOREIGN no04f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 2.985 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.405 0.495 4.240 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.755 0.495 7.690 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 10.125 0.490 11.3100 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.475 0.590 14.310 0.770 ;
        END
    END d
END no04f10
MACRO no04f20
    CLASS CORE ;
    FOREIGN no04f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 33.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 5.930 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.755 0.495 8.425 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.475 0.495 15.145 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 20.205 0.490 22.550 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 26.915 0.590 28.585 0.770 ;
        END
    END d
END no04f20
MACRO no04f40
    CLASS CORE ;
    FOREIGN no04f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 67.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 11.835 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 13.475 0.495 16.810 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 26.915 0.495 30.250 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 40.355 0.490 45.055 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 53.805 0.590 57.140 0.770 ;
        END
    END d
END no04f40
MACRO no04f80
    CLASS CORE ;
    FOREIGN no04f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 134.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.360 23.625 0.900 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 26.915 0.495 33.690 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 53.805 0.495 60.580 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 80.675 0.490 90.065 0.870 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 107.565 0.590 114.240 0.770 ;
        END
    END d
END no04f80
MACRO ao12s01
    CLASS CORE ;
    FOREIGN ao12s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 0.125 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.280 0.495 0.375 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.535 0.495 0.650 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.770 0.590 0.860 0.770 ;
        END
    END c
END ao12s01
MACRO ao12s02
    CLASS CORE ;
    FOREIGN ao12s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 0.2100 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.535 0.495 0.725 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.015 0.495 1.255 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.590 1.695 0.770 ;
        END
    END c
END ao12s02
MACRO ao12s03
    CLASS CORE ;
    FOREIGN ao12s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 0.280 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.770 0.495 1.050 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.495 1.850 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.240 0.590 2.510 0.770 ;
        END
    END c
END ao12s03
MACRO ao12s04
    CLASS CORE ;
    FOREIGN ao12s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 0.365 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.015 0.495 1.390 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.495 2.570 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.985 0.590 3.355 0.770 ;
        END
    END c
END ao12s04
MACRO ao12s06
    CLASS CORE ;
    FOREIGN ao12s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 0.530 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.495 2.070 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.985 0.495 3.780 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.455 0.590 5.005 0.770 ;
        END
    END c
END ao12s06
MACRO ao12s08
    CLASS CORE ;
    FOREIGN ao12s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 0.695 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.495 2.860 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.495 4.890 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.925 0.590 6.645 0.770 ;
        END
    END c
END ao12s08
MACRO ao12s10
    CLASS CORE ;
    FOREIGN ao12s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 1.350 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.495 5.470 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.495 9.735 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 11.795 0.590 13.235 0.770 ;
        END
    END c
END ao12s10
MACRO ao12s20
    CLASS CORE ;
    FOREIGN ao12s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 31.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 2.675 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.495 10.9100 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.495 19.425 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 23.555 0.590 26.435 0.770 ;
        END
    END c
END ao12s20
MACRO ao12s40
    CLASS CORE ;
    FOREIGN ao12s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 62.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 5.3100 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.495 21.740 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 31.395 0.495 38.805 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 47.085 0.590 52.845 0.770 ;
        END
    END c
END ao12s40
MACRO ao12s80
    CLASS CORE ;
    FOREIGN ao12s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 125.440 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 10.560 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 31.395 0.495 43.450 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 62.765 0.495 77.670 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 94.115 0.590 105.645 0.770 ;
        END
    END c
END ao12s80
MACRO ao12m01
    CLASS CORE ;
    FOREIGN ao12m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 0.125 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.280 0.495 0.375 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.535 0.495 0.650 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.770 0.590 0.860 0.770 ;
        END
    END c
END ao12m01
MACRO ao12m02
    CLASS CORE ;
    FOREIGN ao12m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 0.2100 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.535 0.495 0.725 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.015 0.495 1.255 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.590 1.695 0.770 ;
        END
    END c
END ao12m02
MACRO ao12m03
    CLASS CORE ;
    FOREIGN ao12m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 0.280 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.770 0.495 1.050 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.495 1.850 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.240 0.590 2.510 0.770 ;
        END
    END c
END ao12m03
MACRO ao12m04
    CLASS CORE ;
    FOREIGN ao12m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 0.365 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.015 0.495 1.390 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.495 2.570 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.985 0.590 3.355 0.770 ;
        END
    END c
END ao12m04
MACRO ao12m06
    CLASS CORE ;
    FOREIGN ao12m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 0.530 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.495 2.070 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.985 0.495 3.780 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.455 0.590 5.005 0.770 ;
        END
    END c
END ao12m06
MACRO ao12m08
    CLASS CORE ;
    FOREIGN ao12m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 0.695 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.495 2.860 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.495 4.890 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.925 0.590 6.645 0.770 ;
        END
    END c
END ao12m08
MACRO ao12m10
    CLASS CORE ;
    FOREIGN ao12m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 1.350 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.495 5.470 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.495 9.735 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 11.795 0.590 13.235 0.770 ;
        END
    END c
END ao12m10
MACRO ao12m20
    CLASS CORE ;
    FOREIGN ao12m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 31.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 2.675 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.495 10.9100 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.495 19.425 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 23.555 0.590 26.435 0.770 ;
        END
    END c
END ao12m20
MACRO ao12m40
    CLASS CORE ;
    FOREIGN ao12m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 62.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 5.3100 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.495 21.740 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 31.395 0.495 38.805 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 47.085 0.590 52.845 0.770 ;
        END
    END c
END ao12m40
MACRO ao12m80
    CLASS CORE ;
    FOREIGN ao12m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 125.440 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 10.560 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 31.395 0.495 43.450 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 62.765 0.495 77.670 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 94.115 0.590 105.645 0.770 ;
        END
    END c
END ao12m80
MACRO ao12f01
    CLASS CORE ;
    FOREIGN ao12f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 0.125 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.280 0.495 0.375 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.535 0.495 0.650 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.770 0.590 0.860 0.770 ;
        END
    END c
END ao12f01
MACRO ao12f02
    CLASS CORE ;
    FOREIGN ao12f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 0.2100 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.535 0.495 0.725 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.015 0.495 1.255 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.590 1.695 0.770 ;
        END
    END c
END ao12f02
MACRO ao12f03
    CLASS CORE ;
    FOREIGN ao12f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 0.280 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.770 0.495 1.050 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.495 1.850 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.240 0.590 2.510 0.770 ;
        END
    END c
END ao12f03
MACRO ao12f04
    CLASS CORE ;
    FOREIGN ao12f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 0.365 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.015 0.495 1.390 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.495 2.570 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.985 0.590 3.355 0.770 ;
        END
    END c
END ao12f04
MACRO ao12f06
    CLASS CORE ;
    FOREIGN ao12f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 0.530 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.495 2.070 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.985 0.495 3.780 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.455 0.590 5.005 0.770 ;
        END
    END c
END ao12f06
MACRO ao12f08
    CLASS CORE ;
    FOREIGN ao12f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 0.695 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.495 2.860 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.495 4.890 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.925 0.590 6.645 0.770 ;
        END
    END c
END ao12f08
MACRO ao12f10
    CLASS CORE ;
    FOREIGN ao12f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 1.350 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.495 5.470 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.495 9.735 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 11.795 0.590 13.235 0.770 ;
        END
    END c
END ao12f10
MACRO ao12f20
    CLASS CORE ;
    FOREIGN ao12f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 31.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 2.675 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.495 10.9100 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.495 19.425 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 23.555 0.590 26.435 0.770 ;
        END
    END c
END ao12f20
MACRO ao12f40
    CLASS CORE ;
    FOREIGN ao12f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 62.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 5.3100 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.495 21.740 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 31.395 0.495 38.805 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 47.085 0.590 52.845 0.770 ;
        END
    END c
END ao12f40
MACRO ao12f80
    CLASS CORE ;
    FOREIGN ao12f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 125.440 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.205 10.560 1.055 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 31.395 0.495 43.450 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 62.765 0.495 77.670 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 94.115 0.590 105.645 0.770 ;
        END
    END c
END ao12f80
MACRO ao22s01
    CLASS CORE ;
    FOREIGN ao22s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.125 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.295 0.495 0.410 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.540 0.495 0.630 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.790 0.495 0.880 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.590 1.140 0.770 ;
        END
    END d
END ao22s01
MACRO ao22s02
    CLASS CORE ;
    FOREIGN ao22s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.215 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.540 0.495 0.770 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.495 1.235 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.495 1.745 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.590 2.240 0.770 ;
        END
    END d
END ao22s02
MACRO ao22s03
    CLASS CORE ;
    FOREIGN ao22s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.305 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.790 0.495 1.145 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.495 1.825 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.305 0.495 2.585 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.160 0.590 3.445 0.770 ;
        END
    END d
END ao22s03
MACRO ao22s04
    CLASS CORE ;
    FOREIGN ao22s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.405 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.495 1.510 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.495 2.410 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.160 0.495 3.520 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.590 4.465 0.770 ;
        END
    END d
END ao22s04
MACRO ao22s06
    CLASS CORE ;
    FOREIGN ao22s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.575 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.495 2.250 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.160 0.495 3.700 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.570 0.495 5.110 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.085 0.590 6.665 0.770 ;
        END
    END d
END ao22s06
MACRO ao22s08
    CLASS CORE ;
    FOREIGN ao22s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.765 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.495 2.985 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.495 4.795 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.085 0.495 6.805 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.1100 0.590 8.870 0.770 ;
        END
    END d
END ao22s08
MACRO ao22s10
    CLASS CORE ;
    FOREIGN ao22s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 1.485 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.495 5.925 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.1100 0.495 9.550 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 12.130 0.495 13.570 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 16.165 0.590 17.685 0.770 ;
        END
    END d
END ao22s10
MACRO ao22s20
    CLASS CORE ;
    FOREIGN ao22s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 40.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 2.925 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.1100 0.495 11.810 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 16.165 0.495 19.055 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 24.235 0.495 27.115 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 32.290 0.590 35.330 0.770 ;
        END
    END d
END ao22s20
MACRO ao22s40
    CLASS CORE ;
    FOREIGN ao22s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 80.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 5.795 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 16.165 0.495 23.575 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 32.290 0.495 38.050 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 48.420 0.495 54.180 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 64.555 0.590 70.645 0.770 ;
        END
    END d
END ao22s40
MACRO ao22s80
    CLASS CORE ;
    FOREIGN ao22s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 161.280 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 11.555 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 32.290 0.495 47.095 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 64.555 0.495 76.085 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 96.805 0.495 108.335 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 129.160 0.590 141.320 0.770 ;
        END
    END d
END ao22s80
MACRO ao22m01
    CLASS CORE ;
    FOREIGN ao22m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.125 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.295 0.495 0.410 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.540 0.495 0.630 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.790 0.495 0.880 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.590 1.140 0.770 ;
        END
    END d
END ao22m01
MACRO ao22m02
    CLASS CORE ;
    FOREIGN ao22m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.215 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.540 0.495 0.770 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.495 1.235 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.495 1.745 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.590 2.240 0.770 ;
        END
    END d
END ao22m02
MACRO ao22m03
    CLASS CORE ;
    FOREIGN ao22m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.305 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.790 0.495 1.145 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.495 1.825 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.305 0.495 2.585 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.160 0.590 3.445 0.770 ;
        END
    END d
END ao22m03
MACRO ao22m04
    CLASS CORE ;
    FOREIGN ao22m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.405 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.495 1.510 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.495 2.410 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.160 0.495 3.520 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.590 4.465 0.770 ;
        END
    END d
END ao22m04
MACRO ao22m06
    CLASS CORE ;
    FOREIGN ao22m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.575 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.495 2.250 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.160 0.495 3.700 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.570 0.495 5.110 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.085 0.590 6.665 0.770 ;
        END
    END d
END ao22m06
MACRO ao22m08
    CLASS CORE ;
    FOREIGN ao22m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.765 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.495 2.985 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.495 4.795 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.085 0.495 6.805 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.1100 0.590 8.870 0.770 ;
        END
    END d
END ao22m08
MACRO ao22m10
    CLASS CORE ;
    FOREIGN ao22m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 1.485 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.495 5.925 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.1100 0.495 9.550 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 12.130 0.495 13.570 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 16.165 0.590 17.685 0.770 ;
        END
    END d
END ao22m10
MACRO ao22m20
    CLASS CORE ;
    FOREIGN ao22m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 40.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 2.925 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.1100 0.495 11.810 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 16.165 0.495 19.055 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 24.235 0.495 27.115 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 32.290 0.590 35.330 0.770 ;
        END
    END d
END ao22m20
MACRO ao22m40
    CLASS CORE ;
    FOREIGN ao22m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 80.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 5.795 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 16.165 0.495 23.575 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 32.290 0.495 38.050 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 48.420 0.495 54.180 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 64.555 0.590 70.645 0.770 ;
        END
    END d
END ao22m40
MACRO ao22m80
    CLASS CORE ;
    FOREIGN ao22m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 161.280 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 11.555 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 32.290 0.495 47.095 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 64.555 0.495 76.085 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 96.805 0.495 108.335 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 129.160 0.590 141.320 0.770 ;
        END
    END d
END ao22m80
MACRO ao22f01
    CLASS CORE ;
    FOREIGN ao22f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.125 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.295 0.495 0.410 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.540 0.495 0.630 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.790 0.495 0.880 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.590 1.140 0.770 ;
        END
    END d
END ao22f01
MACRO ao22f02
    CLASS CORE ;
    FOREIGN ao22f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.215 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.540 0.495 0.770 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.495 1.235 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.495 1.745 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.590 2.240 0.770 ;
        END
    END d
END ao22f02
MACRO ao22f03
    CLASS CORE ;
    FOREIGN ao22f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.305 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.790 0.495 1.145 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.495 1.825 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.305 0.495 2.585 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.160 0.590 3.445 0.770 ;
        END
    END d
END ao22f03
MACRO ao22f04
    CLASS CORE ;
    FOREIGN ao22f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.405 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.495 1.510 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.495 2.410 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.160 0.495 3.520 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.590 4.465 0.770 ;
        END
    END d
END ao22f04
MACRO ao22f06
    CLASS CORE ;
    FOREIGN ao22f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.575 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.495 2.250 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.160 0.495 3.700 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.570 0.495 5.110 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.085 0.590 6.665 0.770 ;
        END
    END d
END ao22f06
MACRO ao22f08
    CLASS CORE ;
    FOREIGN ao22f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 0.765 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.495 2.985 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.495 4.795 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.085 0.495 6.805 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.1100 0.590 8.870 0.770 ;
        END
    END d
END ao22f08
MACRO ao22f10
    CLASS CORE ;
    FOREIGN ao22f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 1.485 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.495 5.925 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.1100 0.495 9.550 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 12.130 0.495 13.570 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 16.165 0.590 17.685 0.770 ;
        END
    END d
END ao22f10
MACRO ao22f20
    CLASS CORE ;
    FOREIGN ao22f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 40.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 2.925 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.1100 0.495 11.810 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 16.165 0.495 19.055 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 24.235 0.495 27.115 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 32.290 0.590 35.330 0.770 ;
        END
    END d
END ao22f20
MACRO ao22f40
    CLASS CORE ;
    FOREIGN ao22f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 80.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 5.795 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 16.165 0.495 23.575 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 32.290 0.495 38.050 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 48.420 0.495 54.180 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 64.555 0.590 70.645 0.770 ;
        END
    END d
END ao22f40
MACRO ao22f80
    CLASS CORE ;
    FOREIGN ao22f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 161.280 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.200 11.555 1.060 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 32.290 0.495 47.095 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 64.555 0.495 76.085 0.775 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 96.805 0.495 108.335 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 129.160 0.590 141.320 0.770 ;
        END
    END d
END ao22f80
MACRO oa12s01
    CLASS CORE ;
    FOREIGN oa12s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 0.125 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.280 0.495 0.375 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.535 0.590 0.760 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.770 0.425 0.860 0.835 ;
        END
    END c
END oa12s01
MACRO oa12s02
    CLASS CORE ;
    FOREIGN oa12s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 0.215 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.535 0.495 0.725 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.015 0.590 1.260 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.425 1.695 0.835 ;
        END
    END c
END oa12s02
MACRO oa12s03
    CLASS CORE ;
    FOREIGN oa12s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 0.305 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.770 0.495 1.050 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.590 1.875 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.240 0.425 2.510 0.835 ;
        END
    END c
END oa12s03
MACRO oa12s04
    CLASS CORE ;
    FOREIGN oa12s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 0.405 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.015 0.495 1.390 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.590 2.505 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.985 0.425 3.355 0.835 ;
        END
    END c
END oa12s04
MACRO oa12s06
    CLASS CORE ;
    FOREIGN oa12s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 0.575 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.495 2.070 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.985 0.590 3.725 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.455 0.425 5.005 0.835 ;
        END
    END c
END oa12s06
MACRO oa12s08
    CLASS CORE ;
    FOREIGN oa12s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 0.765 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.495 2.860 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.590 4.950 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.925 0.425 6.645 0.835 ;
        END
    END c
END oa12s08
MACRO oa12s10
    CLASS CORE ;
    FOREIGN oa12s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 1.485 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.495 5.470 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.590 9.855 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 11.795 0.425 13.235 0.835 ;
        END
    END c
END oa12s10
MACRO oa12s20
    CLASS CORE ;
    FOREIGN oa12s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 31.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 2.925 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.495 10.9100 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.590 19.655 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 23.555 0.425 26.435 0.835 ;
        END
    END c
END oa12s20
MACRO oa12s40
    CLASS CORE ;
    FOREIGN oa12s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 62.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 5.795 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.495 21.740 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 31.395 0.590 39.270 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 47.085 0.425 52.845 0.835 ;
        END
    END c
END oa12s40
MACRO oa12s80
    CLASS CORE ;
    FOREIGN oa12s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 125.440 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 11.555 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 31.395 0.495 43.450 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 62.765 0.590 78.520 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 94.115 0.425 105.645 0.835 ;
        END
    END c
END oa12s80
MACRO oa12m01
    CLASS CORE ;
    FOREIGN oa12m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 0.125 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.280 0.495 0.375 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.535 0.590 0.760 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.770 0.425 0.860 0.835 ;
        END
    END c
END oa12m01
MACRO oa12m02
    CLASS CORE ;
    FOREIGN oa12m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 0.215 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.535 0.495 0.725 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.015 0.590 1.260 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.425 1.695 0.835 ;
        END
    END c
END oa12m02
MACRO oa12m03
    CLASS CORE ;
    FOREIGN oa12m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 0.305 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.770 0.495 1.050 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.590 1.875 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.240 0.425 2.510 0.835 ;
        END
    END c
END oa12m03
MACRO oa12m04
    CLASS CORE ;
    FOREIGN oa12m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 0.405 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.015 0.495 1.390 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.590 2.505 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.985 0.425 3.355 0.835 ;
        END
    END c
END oa12m04
MACRO oa12m06
    CLASS CORE ;
    FOREIGN oa12m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 0.575 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.495 2.070 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.985 0.590 3.725 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.455 0.425 5.005 0.835 ;
        END
    END c
END oa12m06
MACRO oa12m08
    CLASS CORE ;
    FOREIGN oa12m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 0.765 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.495 2.860 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.590 4.950 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.925 0.425 6.645 0.835 ;
        END
    END c
END oa12m08
MACRO oa12m10
    CLASS CORE ;
    FOREIGN oa12m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 1.485 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.495 5.470 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.590 9.855 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 11.795 0.425 13.235 0.835 ;
        END
    END c
END oa12m10
MACRO oa12m20
    CLASS CORE ;
    FOREIGN oa12m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 31.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 2.925 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.495 10.9100 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.590 19.655 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 23.555 0.425 26.435 0.835 ;
        END
    END c
END oa12m20
MACRO oa12m40
    CLASS CORE ;
    FOREIGN oa12m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 62.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 5.795 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.495 21.740 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 31.395 0.590 39.270 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 47.085 0.425 52.845 0.835 ;
        END
    END c
END oa12m40
MACRO oa12m80
    CLASS CORE ;
    FOREIGN oa12m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 125.440 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 11.555 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 31.395 0.495 43.450 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 62.765 0.590 78.520 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 94.115 0.425 105.645 0.835 ;
        END
    END c
END oa12m80
MACRO oa12f01
    CLASS CORE ;
    FOREIGN oa12f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 0.125 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.280 0.495 0.375 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.535 0.590 0.760 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.770 0.425 0.860 0.835 ;
        END
    END c
END oa12f01
MACRO oa12f02
    CLASS CORE ;
    FOREIGN oa12f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 0.215 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.535 0.495 0.725 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.015 0.590 1.260 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.425 1.695 0.835 ;
        END
    END c
END oa12f02
MACRO oa12f03
    CLASS CORE ;
    FOREIGN oa12f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 0.305 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.770 0.495 1.050 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.590 1.875 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.240 0.425 2.510 0.835 ;
        END
    END c
END oa12f03
MACRO oa12f04
    CLASS CORE ;
    FOREIGN oa12f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 0.405 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.015 0.495 1.390 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.590 2.505 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.985 0.425 3.355 0.835 ;
        END
    END c
END oa12f04
MACRO oa12f06
    CLASS CORE ;
    FOREIGN oa12f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 0.575 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.505 0.495 2.070 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.985 0.590 3.725 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.455 0.425 5.005 0.835 ;
        END
    END c
END oa12f06
MACRO oa12f08
    CLASS CORE ;
    FOREIGN oa12f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 0.765 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.005 0.495 2.860 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.590 4.950 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 5.925 0.425 6.645 0.835 ;
        END
    END c
END oa12f08
MACRO oa12f10
    CLASS CORE ;
    FOREIGN oa12f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 1.485 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.965 0.495 5.470 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.590 9.855 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 11.795 0.425 13.235 0.835 ;
        END
    END c
END oa12f10
MACRO oa12f20
    CLASS CORE ;
    FOREIGN oa12f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 31.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 2.925 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 7.885 0.495 10.9100 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.590 19.655 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 23.555 0.425 26.435 0.835 ;
        END
    END c
END oa12f20
MACRO oa12f40
    CLASS CORE ;
    FOREIGN oa12f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 62.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 5.795 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 15.715 0.495 21.740 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 31.395 0.590 39.270 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 47.085 0.425 52.845 0.835 ;
        END
    END c
END oa12f40
MACRO oa12f80
    CLASS CORE ;
    FOREIGN oa12f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 125.440 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 11.555 1.070 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 31.395 0.495 43.450 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 62.765 0.590 78.520 0.770 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 94.115 0.425 105.645 0.835 ;
        END
    END c
END oa12f80
MACRO oa22s01
    CLASS CORE ;
    FOREIGN oa22s01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 0.125 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.295 0.495 0.410 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.540 0.425 0.630 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.790 0.495 0.880 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.495 1.140 0.775 ;
        END
    END d
END oa22s01
MACRO oa22s02
    CLASS CORE ;
    FOREIGN oa22s02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 0.215 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.540 0.495 0.770 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.425 1.235 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.495 1.745 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.495 2.240 0.775 ;
        END
    END d
END oa22s02
MACRO oa22s03
    CLASS CORE ;
    FOREIGN oa22s03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 0.305 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.790 0.495 1.145 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.425 1.825 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.305 0.495 2.585 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.160 0.495 3.445 0.775 ;
        END
    END d
END oa22s03
MACRO oa22s04
    CLASS CORE ;
    FOREIGN oa22s04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 0.405 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.495 1.510 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.425 2.410 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.160 0.495 3.520 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.495 4.465 0.775 ;
        END
    END d
END oa22s04
MACRO oa22s06
    CLASS CORE ;
    FOREIGN oa22s06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 0.575 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.495 2.250 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.160 0.425 3.700 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.570 0.495 5.110 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.085 0.495 6.665 0.775 ;
        END
    END d
END oa22s06
MACRO oa22s08
    CLASS CORE ;
    FOREIGN oa22s08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 0.765 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.495 2.985 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.425 4.795 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.085 0.495 6.805 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.1100 0.495 8.870 0.775 ;
        END
    END d
END oa22s08
MACRO oa22s10
    CLASS CORE ;
    FOREIGN oa22s10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 1.485 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.495 5.925 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.1100 0.425 9.550 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 12.130 0.495 13.570 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 16.165 0.495 17.685 0.775 ;
        END
    END d
END oa22s10
MACRO oa22s20
    CLASS CORE ;
    FOREIGN oa22s20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 40.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 2.925 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.1100 0.495 11.810 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 16.165 0.425 19.055 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 24.235 0.495 27.115 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 32.290 0.495 35.330 0.775 ;
        END
    END d
END oa22s20
MACRO oa22s40
    CLASS CORE ;
    FOREIGN oa22s40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 80.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 5.795 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 16.165 0.495 23.575 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 32.290 0.425 38.050 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 48.420 0.495 54.180 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 64.555 0.495 70.645 0.775 ;
        END
    END d
END oa22s40
MACRO oa22s80
    CLASS CORE ;
    FOREIGN oa22s80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 161.280 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 11.555 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 32.290 0.495 47.095 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 64.555 0.425 76.085 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 96.805 0.495 108.335 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 129.160 0.495 141.320 0.775 ;
        END
    END d
END oa22s80
MACRO oa22m01
    CLASS CORE ;
    FOREIGN oa22m01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 0.125 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.295 0.495 0.410 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.540 0.425 0.630 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.790 0.495 0.880 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.495 1.140 0.775 ;
        END
    END d
END oa22m01
MACRO oa22m02
    CLASS CORE ;
    FOREIGN oa22m02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 0.215 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.540 0.495 0.770 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.425 1.235 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.495 1.745 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.495 2.240 0.775 ;
        END
    END d
END oa22m02
MACRO oa22m03
    CLASS CORE ;
    FOREIGN oa22m03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 0.305 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.790 0.495 1.145 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.425 1.825 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.305 0.495 2.585 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.160 0.495 3.445 0.775 ;
        END
    END d
END oa22m03
MACRO oa22m04
    CLASS CORE ;
    FOREIGN oa22m04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 0.405 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.495 1.510 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.425 2.410 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.160 0.495 3.520 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.495 4.465 0.775 ;
        END
    END d
END oa22m04
MACRO oa22m06
    CLASS CORE ;
    FOREIGN oa22m06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 0.575 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.495 2.250 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.160 0.425 3.700 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.570 0.495 5.110 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.085 0.495 6.665 0.775 ;
        END
    END d
END oa22m06
MACRO oa22m08
    CLASS CORE ;
    FOREIGN oa22m08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 0.765 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.495 2.985 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.425 4.795 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.085 0.495 6.805 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.1100 0.495 8.870 0.775 ;
        END
    END d
END oa22m08
MACRO oa22m10
    CLASS CORE ;
    FOREIGN oa22m10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 1.485 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.495 5.925 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.1100 0.425 9.550 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 12.130 0.495 13.570 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 16.165 0.495 17.685 0.775 ;
        END
    END d
END oa22m10
MACRO oa22m20
    CLASS CORE ;
    FOREIGN oa22m20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 40.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 2.925 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.1100 0.495 11.810 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 16.165 0.425 19.055 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 24.235 0.495 27.115 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 32.290 0.495 35.330 0.775 ;
        END
    END d
END oa22m20
MACRO oa22m40
    CLASS CORE ;
    FOREIGN oa22m40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 80.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 5.795 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 16.165 0.495 23.575 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 32.290 0.425 38.050 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 48.420 0.495 54.180 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 64.555 0.495 70.645 0.775 ;
        END
    END d
END oa22m40
MACRO oa22m80
    CLASS CORE ;
    FOREIGN oa22m80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 161.280 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 11.555 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 32.290 0.495 47.095 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 64.555 0.425 76.085 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 96.805 0.495 108.335 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 129.160 0.495 141.320 0.775 ;
        END
    END d
END oa22m80
MACRO oa22f01
    CLASS CORE ;
    FOREIGN oa22f01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 0.125 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.295 0.495 0.410 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.540 0.425 0.630 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.790 0.495 0.880 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.495 1.140 0.775 ;
        END
    END d
END oa22f01
MACRO oa22f02
    CLASS CORE ;
    FOREIGN oa22f02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 0.215 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.540 0.495 0.770 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.425 1.235 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.495 1.745 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.495 2.240 0.775 ;
        END
    END d
END oa22f02
MACRO oa22f03
    CLASS CORE ;
    FOREIGN oa22f03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 0.305 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 0.790 0.495 1.145 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.425 1.825 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.305 0.495 2.585 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.160 0.495 3.445 0.775 ;
        END
    END d
END oa22f03
MACRO oa22f04
    CLASS CORE ;
    FOREIGN oa22f04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 0.405 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.045 0.495 1.510 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.425 2.410 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.160 0.495 3.520 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.495 4.465 0.775 ;
        END
    END d
END oa22f04
MACRO oa22f06
    CLASS CORE ;
    FOREIGN oa22f06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 0.575 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.555 0.495 2.250 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 3.160 0.425 3.700 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.570 0.495 5.110 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.085 0.495 6.665 0.775 ;
        END
    END d
END oa22f06
MACRO oa22f08
    CLASS CORE ;
    FOREIGN oa22f08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 0.765 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.050 0.495 2.985 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.425 4.795 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 6.085 0.495 6.805 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.1100 0.495 8.870 0.775 ;
        END
    END d
END oa22f08
MACRO oa22f10
    CLASS CORE ;
    FOREIGN oa22f10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 1.485 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 4.075 0.495 5.925 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.1100 0.425 9.550 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 12.130 0.495 13.570 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 16.165 0.495 17.685 0.775 ;
        END
    END d
END oa22f10
MACRO oa22f20
    CLASS CORE ;
    FOREIGN oa22f20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 40.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 2.925 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 8.1100 0.495 11.810 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 16.165 0.425 19.055 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 24.235 0.495 27.115 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 32.290 0.495 35.330 0.775 ;
        END
    END d
END oa22f20
MACRO oa22f40
    CLASS CORE ;
    FOREIGN oa22f40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 80.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 5.795 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 16.165 0.495 23.575 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 32.290 0.425 38.050 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 48.420 0.495 54.180 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 64.555 0.495 70.645 0.775 ;
        END
    END d
END oa22f40
MACRO oa22f80
    CLASS CORE ;
    FOREIGN oa22f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 161.280 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.185 11.555 1.075 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 32.290 0.495 47.095 0.775 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 64.555 0.425 76.085 0.835 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 96.805 0.495 108.335 0.775 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 129.160 0.495 141.320 0.775 ;
        END
    END d
END oa22f80
MACRO ms00f80
    CLASS CORE ;
    FOREIGN ms00f80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT 0.035 0.190 0.290 1.070 ;
        END
    END o
    PIN ck
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 1.445 0.495 1.535 0.775 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT 2.835 0.490 2.950 0.770 ;
        END
    END d
END ms00f80
END LIBRARY
